XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����٬�����siO"i�&P?<�;�ߨ��a�7��s��9��o�,\ӓC�2Ve��#'�[&���T_#���8��.p
xW��_�U䋩2�u�.��.!��0н��� p�z��� ��7�Gr���,F����� rG�D8����6-����f ��ł��m]���gF[av���N�ކ�����&�ڻK�4�^zU4��R�V M���mR���!@�m�Q��y+�:Y���S�"��Pu&����I�l�/�u���
�&���t!X��P]gm��M.��ˀ�|�O��.�'p�^j��l@6��&���jUȜ�yA���%�ݴ.vA��E�g�>���Dp2�����sf��!�T��K��zd��ŀ~���(uշ��xͬz�Lגn#��e[?��2q�`|HU�K����a�2^6�)?���>�2_Zv��R���y]X�_?>o�N��"����	X.lY&7�`�O������k�H�w�$y�%��i�R�>�`޺Tև�/H������`�M�(��� b��K�э�T)>���E\i���b|��B���Ħe���S=T��#$���=��ʹ[]5�+�6ޔ��:���!�Ě�Z��#�6]�euS�%�NV�����uk�̼�����;��ȝͼ�
�_7t����"/y�/�u�_���6�8�	�N��v�|����+���ޛ&���!����tB��L^y�09�����/�F�YG�����XlxVHYEB    5b61    1040��1�+%�Zԇ���쒅+@��Pn:7v!�GN�W$�9e_���fu!�F��%�(E�W�,v_��n��_y2�$���0�Y��A������&>�`��� �5��9����{�,�k���/R/�g0�Gڬ�����t��7,%��W��|^���d��W�����L��*�\#U���س1 w-�ȝtu_U�nߒݯgΕ��j^XZH�����"%���`�����/h����k�k��F؍�6��]�7�SwP�P��8;<�E9�0tO&�'�,�L�}kx���)֮MK{�jަ�`%Yn�~�<�'=,�Z�z��@k�:U��u����0>�(���-��s��M�4ݡ6<?���JR��,�; �bM^���`�ES-�n:�DIiukW'��b����[����{��������˗:}�f[S�S5_m��7	��j����d$�}�iRA�� ?�k3��=	,O*K4~��F)r�U��\k���ι�
L��I�y�W���x�{&eX���0�u��=c��B������1�����Lqϝ�}w�-
�����	�3��h ��C���gz�a�8K�d���'�Rj�;.�������V�~9S씣��Tg<��N3��m������!��ʉ%ʔk���i,I�;��f�Z嗦8�BF?mNS����l�(yk��U^�����w�+ s��6�~���Nd�D8.������*�C��l�/���6�6c9��*�\�!�A	���5��<���Vb�kʼu��"�7�3X˦�MOr��ܶ���0�7Ν:��Ϥ�����N�*���B\�]?m=L�rh�7�庢��a~����^���#��h�^��g���Poa��紹��G����*�_y�	����$�sg�w�bW�t���ŗ�L����|&q��ʜ���O]��XY5a����liwHE�����0���y�s6���ԗy�7�>�dz:IE��\��S����\0����-�*� �v��RM��B�l��(F����Ʒi5ɼr&��G����X��}c�g����-ַ�DD��\p/X�3�)gK}��fɹ�4�Sl��s}���U?�]!�`���Ϊ$䊩�Ț�$s�o�ȼ�
�BB�A���H  _������Q�!2{HK��\�V�gh=q3'�sH7j'�&u�,���f��@�cr_��/�\�y3��@4�:�=��!��`�k��=l#K��~�p�?��N�'�S��!�P6�v/'�~F������gz�����Lk�9D&aʇ��`�Q��_E�O\'�	���S�M<�IGA�5֗�!K�@�#����{�j*vR�M��%�_�/�M��FΟ��/�AE���W�'�"F)����\��3���g+C=�#1�֝�^�/շ�p=kh�����i(��O�ڈ����p�Rő���»�Ļ�01�Ӆ�V��<���cġ�塴�;�N�zW$�?�&v�n���(�����.��.՘�����C�w��{>���� v-�"���f��l_�	�"=�f���I�,�5
�H8֮}������BuA��ܢn���}�L�¸Ml�;cF���jr6�H&�G�?hI�?�@�h�#5�*�z[�+�F���u������h����;^���z��w@���neu>����B�5b�.��n,$'6��_P���5�U#�2�����#w�h�y+���u�ސK���c�Y����J�A�r�.໲���e�g�,�m(�R���X���X�*�S�* 39�A�(���|E�@���nU�8�(H���2��yHQl�}���������{���{�֋�ד����w�BL�@��
>1[\�Y�e@7��V�I%�޾�\�D��)g��aY��ȑ??�a%=?X�r�͌��S��rs���,��Uϔ��IQ�'��+ܰ.��,�b����Ce���@��_��{��f��PI��}5��:�I������5Kh��:;G���2!�Q��[�OL%Vy�_fM/�G9v��˽Y�M���oߓ8�GIe��yq7 V,�4"1�
��0�3*���3���ؤF�|@_���ju��=6�QI�;�e��<M|��8m���y!��$JN0�LҋX�9�����No�}K��r���R���_��6��a ���c���{��Ț�B���e�^ʲz��M~_����I}M�ksx=� n��h��~�a�%v�������ԛ�$��Q��x���$�0�E�_ƲU#s����@��P���k1��dq��"Y4�.g�Xy��`��^��,�X
 ��6�1c�C�����,�ݛPFW5-F�o�W�]_�a�PV�0w�f2�H3���W���N���`����
����DI�t��I�⼏�HD\��Kj͕���W�6�=�N��`�����iI��cI��Y>9�EDޏ �*�_t~\� (�O���2�����]��k�4u$�"�
G��nPR-���|��=2�/`U�Äb�jzԬO�Js犋Ż}�B��#_u,�$����������,>ي8���؝�P���]�����Wfq7�� !]�q���n�)qe��i���?M&)`��D:g���g��;����1���� �g�>��1Q+�ݹU['Դ�w���c޻rP�1=T��o=W��q3fV�L��$q��W���v��7�t�ga�w�6c���HW^X}��  �#O���{���q�+W�^��l绱d���.�Y��2�?�kgezR_�x�)s{o'�9k����	P�����'�kc�B?_iN��*������0$���E��U�!����]U�=��{X⥞Iػ��W;�5FצCQ <;��'����.�NOhocJ���R�%� b��[�@�]��'�x��_�n���= �63c�9��� ��Hͥ�f�R��^��C���)��û9f�J07��|j\�L���0���z��P�-�M4�{�P\�n����Gh��)%Lkc6�d˦~�\Y9�U���sB��A6Saj�{cI&��WZ��N#l��Y�!����J��<�O���۰� �����6��<`S�ÇJ�(adN�0H��-���(Y��?_�e�g>�t;vS.[]oM���WoK�ԥ���ʰ�a��b�x~�1&�މ��r�C3�c��K_��9n����ϐ�H�ұ@��6H�e��`�ǃ� )�àAZw��\�ฃmW��eoB+~�"U ��!p�f�§�qw�� �=��}s�3�5���������0���`�q��	���z�N��Ÿ���F)W�k&�Qp�z+���
	�`�J�3f+b�W������A��C����
��l+�`1�pq�JvY�Pk���/��h@I����m�1Բ1L&"Ҋ=�Mc���H&k��A@��;�;�:D�V���^B�hF�j�&�C�F9`AX�����0Vx��͒f�T�l�d�p�㯑gR�g�%��	�sD�X@��*��	�OHA+�Og� �e�{�1��.ۋB7'�����x�/�K	\�^Y��˃96c��s���[E>,$�Hn��
3�'ZrRދcp��q����
d�j-=~�&&�%P}�[��#��p�P� 2RCg��3����i,CƩ~�t�� wN �j�&�6D4�3�4�Ԏv&j�u/h�ɏ��I��3���ah����e���5BtUa��j��4�i�g7�rzqY�UW.���.Z�����_�����w����9���KR<�P��tJU�u)��v�R�o0K.'pvB l�F-��o����Q&�}�;5,$	��Y]���?~)�_6��ku� 3{"��7��M+�R�m������c��M��ݬ���-~H*l��$`i��5�p8^����9{0 .�|��|{��	2p��Z��}�+{�iN�w����K/�V=Ӕ��":����cF��������I˚���$�5��׎o��R��U 
��l ^����U��ښ<pbUg_�	�i��*���r��\�v�l��{�� d/WS�U�|�K#5�\��p�8I��#��