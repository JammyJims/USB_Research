XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-���~mv��[�a/�p�I+�C@{ ��TUȀ�ߐ���C ^�*{����,:/�_��N��/�1Cz�� /�¯�&�������)��W�ѱy��|���=~m��|<ԭ$�_#��'3�0W���$�R�I�����7�yb��y	<�b�r`��d��2,%z�٬j���da ���쒤��U����$Ʌ�}q3����e�!��_zB馇��Ϟ#�vԣ�0����Q�)Ë��Vw� *��O�/�?���R�0u��i����xG��4��*^y���,5�ʍ<�rKOK0h�r���#[�e�=�j����ٔ7�/�ޱj{W�9���y>@M�@F<v�q��9�����j�t1��V�v%�ԏ�ȴ-���_��l��,cXs���t/����@��0åg(&�WB g|�z�z0@P9�X獛�=f����	���8
�n���67-5��5�uk���Q�;݉^�K�4U ��>Fz牏��_5ȨTlL?8�Ø�,����'@:zo��o�,�#�)"HԱ���ı��ʄM6�΄;�D���&�ʘ��}�hFI��ڈ�XG2!9��'=��hd��˟�:'� OnW�pӕF±z̩�v��btH��Y�MԬ Ϭf~˾���=g�	QI�I���'�(��tB��K��X���|�.������S����+������!�����ı�Ln.7@��gT����mܚN���a�'�"�F	*8��i�d�6�)�G9O	�'uXlxVHYEB    32ec     940ߩf�����~��d�q�ok��p�����;>$�ݺ�$L�+«���<��; ���u�l}����@
oi��F�\D7�i�j:CJ�m�]O�#7��&vi�W=>w� �o����,��zZx�CD��|W�vŧ.������>*U�x_��~�j�f�JK��82� t0�����FJ1b�cЧKE��Yj!�2�@g��˪0�*DZ�Љ�A#x(ύ%�i��X�ԽY�)���ۑB8|��S�>��9�?o2�am�1�(oq�)C�Ȏ['�^��[	��2��Ѕ�sK�_�_��1��(_=AX�.eh�iq'���q�;s,��Y�����З߳f=�p'FO�}��x�ئh�Տi*Y)[c_��J�i�s�$�7��f�$������Kș��|��˘�� ��X���/���)�|w�q{�N~�z���1��)sY�"�cp�r�K`ff�\U�JG~KJ�'��;+۟fǦ�z�>�ۮ��NwH	t��c�q����<m�9�
�(v<90Xbiz�ё�i�,�?zà2&X�a'������D�����y��zs�<�&@W>��@�r���֤(�ʬG�Ŋ��ǐ��ٝ�R]�{4��(���
��(k������Bw�`�K\-Wٱ=������ud�'C�G2�`3����Ε.�?BɌ�ezp�[���@)갾�T�j���m^2���V�y��
����]�.��\S����;L��?3< ��G���ah���Vd�M�E%O��6A[A��8�čMU��u��yS��G��a��P5�~^�/1����o�u������\�~�޼��:������I�j�L\�c��-Si�qI���{��d'�]� $T�0D���i�������(}1o�><kШ���:!�i-;��jcx�!+
��+o��z�+��&��nd��mL�3ta,z(�;˗|���-�p�v�t^���p�ʃ �)[5�
W����{����AKfc&�T,�ћ�9�R���R��&�}�/`�`��[��bC$������BgΨ�1�3 �q-�Q�Z�H�w����5�C�8�8@3�W1o��&� tf��S ^����@!�3߷6q1��h�����w3vx��5�TK�MvU�x� ��F@�N昭ɇ�Q/ʑv��3�=z;���`��qT�<y��C��٩�Ȩf�yS1�h�m�e�uϩk`�������OB��{{光�m��zf���56`��r��d��|d>9s_���B�^
w�-�D�ŷ5ʌD�:o�^�v)�Է-ۖ���5`����ȟ��h,C�ܛh����b����c�;9�-�7�j윯{�M^��4!'B�?�A$-���X@U��%e�����E��ḵ�z]ˎS�����,lʱ��;~d5?g�㈿�����FuC�^厱�X$�
�ܿ�*��;�.�"��_�rZ���������(k�0�� ��^4_T:�m'�@�݉CB}�
��p���V}�ߔ��O�~ow��_�Q����Y�#b�e3h_�XR^��3)�zp��t���O�S!��뭼^�̼UYрc�$ů�کH���]�f��O�o�K����Lz8�y�/�	���)Y� �*�}4������J�R�M�V�N�"ح,%�$:t8�ҳq��:��*HO��<h6!�a�=-���/�,OQ/#�<5A�2��ónJ�:˶N6�C��E����Q����zOstnhfWЪSn_$�_"}f.����k�.�O%ie�K`����1O�ebC�ݔ�'W��y�q��,�&#Or�����=}�]��s�B��w�c����Qb�
�=.Q����=�RP�ף�ȭy��KPvS��!eUlr�`�O�/ѼZz#Ӹ/�cr%"�r��.�����c�����2��Ebe�^���`��9��jE׍U��z PUr�`�w��́O1��r��*��Mfp��p~�ϳ�<|�Yݙv��8>��A6nV�6�~���������O�A��(qm�ڙ��=<13�Ki��ɺ��u4��
^�G������0R���1��Woh�^ׂLN�\�?7�����<C?@%�䈕d�U�#�雦��u�[���*��V)�Sx���I!
i���<r�Q�V�
 ��ӱTs3学�b���f��%��E2Y�)�n����A&�z��/�r����c2��|`�*%�V�m�4��Eō���>����a�]E�3�^�Y羌d�ћ�w�b|8u�	_y�j@?�\9��bpra@Q�����M ����dR�H:`�c)5�p�
%p�TS��hjvo�ߧ��凘m�