XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X�D{-��3�J�5`�CQ����^��A3�lǔ�[�E\$d�E
;�Kw�X��aB��E,�:#�-�-���>��zܽjކWh`����j���
� ]��`-�� 8��y�Ph8E��ls!"��!ui7��Qӝ��`�?Ǯ�a����x�$w@?��z��B����Ĳ{C�{�C����a�I�9�B�Ta����[Ql�Hԉ#�R@ �u��{�@O����s��X�t��\������ѿ��-c��a5�D[~rP�煑ʑ�SZ�w���,:�	��Ǯ+xŗ�_z��9gwo 
 6��-u�bm�,M%}s���-�`� �^�p�ĴS0�kɵ�J=v%�����Mh� ����d�s�M�`�N7�8��.:�﮵�~�� -6hͽ�*o����Wk���Q�*��,B��h^� �L���3����!��ޢ�e�^_���W�rbN��..�}�ۜb`����<��tN)�,�2u��DǓ@�������̏Ԡw�#��IE����^v�һ^�m�F��H�sr5����/*��A��e�B��ޭtU�lNz��־��a�m��9�)#N���m7�|-��3bT�w�����{)�Our���+�c<n���[u�	
�4Zz���h�h1��pAOō��w�d�J�вq8�,3��·�}��(�[�Di�7������o��S�+�eI��,��'h���#�ui��p r��X���ʴXE��p���)|��,O�E�pf���t�l+�ݯ
R9��XlxVHYEB     a68     2e0cP�iLF���oe��ǸF�X��oI�w7»��Lk¦Mp���c��f���j�p%��N:�&(��ii�B�X$��m��ڔ,�r��r��"�F>���&i���+�<�2��T��.<ʗ��f�I��N�$C��^q�Bk�czf��T�F�Ԙ��q�55tG��-�����7��w��_�"�&���%T�tz��Ă����T���}rK!�SI)�@0U�7�Ƕ�Qt5PkV負�׸ �X�d5@u�&1,u �����,� p�҆�p���n�y�q���ѿ��LG�v{��1��l�l�[W�h��� ���2=�ANE��*0�=�B�K� ��<��y�����s��E8�U2�����ow��Zn#��}�Z�����#���ݧ�F ?����A\���0���ɱд��l����0'���TUЅh^�����3p'ڶ���/swHȏ&�?IӔ.�X:Ԏ�>�1s̃p�cI-�n��qp�T��.gQ]������v��$2?�O\&Ox�}���?�z�؊��h|w��A��c�޴#̻4d�q��	�{��ب,�B�A��%��-��Q�c���!�Z+_y9�'>�~$c�or��yg%=m�Pp�[s������{�yL��kI�p�ڧ~}�� Q� tǧk&����IG�U���s���ggz3��/�_��
oK?kی�c⊦�8��s� ;�DCYm��x��_6��9�