XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������Z'"*��1Z�9)��4)H�&ЃA�����;[k@m`Dѫo�&óB�����Q�� ��Ǡ�1@s�a�<!>�D��>��w�/EGH���C~\�V��qmJ��(�4��[V9���kg�]�uq.��k�N�uI�?y�fSs�>�ghF�۠*J3�h�y�\������(�w�FWc��k�^����L!�]���p�ȶ�M$�>�{c�$����g��"$�I?]OŐ&��rjW۟q�i6ZP�hE�&��0Y=��'��k�#�N�H����Mud�&�c��w/je��?��X;y�2���l����X�C�
(�3�P^V��b��Mˎ'��Zу���v����ۥ����W~I$�z��|�^� ���0�C���1��E6Z��y��cQ_9��j\�Q$P �&	�a�TQ�M��8VrB��Y��y�׈�q���Sf��Ұ����\��/4�"�+���en�$Lh�o�]o�頋I0���0��}�B��~o4���C�ov���W���SWЪ:�|h�^�ѪY�n��L���ׇ��7	х�B��N4"o�ۑݳ����6G�<��
G�;|��T֢������4��۩Ee>_Ѱ�fz����%A/�����tg`���hqE߸��-���8���|]/H���������dŰ��'��������Kʶ�B߷����~E��6��uF����x��pjQ��B+�i�x~߹r�r+ZB�c��˄�TQXlxVHYEB    938c    1610{��;�������j��a�/ 
�� e�÷�
纺�[M�ߔ��S:9���*��^D�4��SEō��	���&SF�4OEW6_��rwYR�s��A$8�r��g�7I��`�)���j�6� �;z>���W�T1�'�J��U�R?0�E�N@5�
B��r���Z-GQ��.��H@+�,r4Z���U��L�� Xr�9��#��+�}�u"���	3N���F��i���v5h �c��4(��>�|?��V���?&Z2���
���{�!L�/�����:�5>咞�@��щ"!CǨ�1./��9/%m)�K��b�cX����ri0�Tyԁ+�r+�M�E�R������(|W�o������%8k�t����<�=��!!p$⢙��n#��f�7�X��{��y*OGh!YRjf���"��q�����F�D���:�m�)aE8M�f
�x��l�����&�HRKk�>_�����(�T<O�76a�Z�bg�N�"�d��y�9����0��D�9�4̅�~��H������O-��Eq����"�ԣ2�T<�[�0�v��B��>X�C�K�T�@�)����Rq���f�9��y1��q�D�kL�(B`Rh �N�����S�`�T~W�
�=Ft ��
�U��|L��Ռ)7d�"Һ�1��i��]�׳w�3Xĉ�C�0t��ߤ����ۛ+D�<��ty�X�C������E>���.ߩ�;�Me��a�X��ӛH��7"��!,��q� �͍(U����0��x��3����VD�4��󴮔E<�}c���=ͱ�\%Dі+��.�&Q$ܠo����g�bl˧J�E@r?n�o������p�[�*1������z���
�md!]��V�f��=`2@N�!�Y^�s]aub�3SY-�M���� ]�� v{��^u�ۤ�(�Q��qnCD\�̤S-!�у*Vw/�:���Ϯ�y�Lnv�y##zk�i��&O��7��|�F\��J�tt,*�
��fkq���˻����v�p�)�����\��s.CF��7to�ٗ-�+$���0�b7����a�!�$})���%8�0�k��r߹7Ӌ�>Y!s �pq���o�C/ٳA.i����=J��G�(b<*���deX�W� g�����t�[6����� _��51��+l)X����M�2.�M��ǳf�m7���Bu\s�me�`�b��|�P=%#o#am.(b?�;¿�v'��B��\�ܼ��Z/��8���M���J���ȴ[��	g�tz�A�����klE �.�������"�!���b��0"Z�a��F�(������fl!Ϗ3��n�T��U$
Q�S9����Y��B�ɡ���u���Z�y�����OM��0��n0>�F�l�%�.���Ȇ�:��Q��e:d���}���*<,�����*/ە�0/�o<vI�q�Is5����-)Kq��t��31�Rz^T&�f�i���\��j��
A�{��"�h�[q)��@��[�d�g��V+�\
L��V���dŎY�܎���!Ԥ����.��Lؚ���!^,J>bEc"�L���5��V��q���km</o�Ƒ�UW�tS	/�6��{%�-kF�=�HI�~B��Wй��E�k�	�w�F�<�ex;G���#�o)[d��ݏ�+��і��5  l͇�׊�/DX���f�h�5�L���ne @n����/��	9�i��v�*}{��)�5�P����=��"�	ˠNh�+��p*E*��b`�!hF}G�N��X��X(�[�-k!��'~)�*��(����[Z�s!�9[pA��x�y�_�5��)����.!��E���*��	���7��hҚڔح+�/@#U��Dz{{@8��%hj��w�Z���z=�;�N�E I. >�	���Ɉ�j1��C��m0��zLl�������� ��H5�lJ�7ԃ\#��Ӷ�
�����T�he5�n���#�Xp��DÛx�8X����n4Nt�m�k���5��������.�M��Sn�$�q�t�%��f����Y� ڷ����f�������PU������m�E·QP]8U)K��Nw�АxIF��&)$��[^�މN/���A��|W)�z "{�xݱ���k�jn[�c��Mb�'0�M5��@Kf������Ȫg<s9<L�� nr��+�~��D</���n�f�м%�į����������K�����s$r�w7ER:a�L���Gg����Uc*�B]̞�����	�+>�%XϰS�h���R���~ß�s}��yքٞU���C'�v}8X�Yg-P�)7Ի�_�؅H�:���m�̭7]#�0ԝ�cH_��;�4K�ۛ�:��^��jV^U��� ��]�C��u�H��t�����0FR�
2MZ~R�{�|��Ջ�U���վҹ�L"�����ҍ�/k��JX$�h��P_��Uh����g�E/ٜUc�|���!���yh���C��P��'��R�3Fm��[fs{���,�Hj��p�۠�w`�y�C)Ds  ��Vl��EG���q��[�TF�_�{�
LB�� qC&��^X�++¨a L7z��qZ�o�	W�"kى�(!�aOѡ��3��sL��o�u��W�fJ�f�0C�p��8T�1�x]��<�KYc�'���̌Z�i�o�_���ٗX�'>�׼��܃RDy�n���5�>��t$�����hJ+���.rj��}"���ͣ��Wt��_�����u��N�4>�`��?/IY���\ҽ����-����x�j����|1���8�ԟW*m�����*�I#��d>0�D��V~`��Ė�j���*�*e�K�}1���Z�v>�v�/��0s(|�:[ S�H^"�}�Uy��ު���d%tI���h���>R��j�2����@� ����I����x����e�k��c�Z�Z��_��A,<=�ъ��<+�6�ˆ�ƥ�S�giQ�����`�N�5�7a�!�}��a_J���b+.��ԑ-�7�1gB�;�?)�n��e@���۶V�_�C�](����=�!�?&��σ�[�����(h�� E_��ɫ��$�|^�ܖ�(\bu���'oD�6IK���B�@ygq��u���ٔ�D��Z*�{�"��z��Uq=#7O:2�b�GKkA
�g�@� (o�7���RUJ;�o5�BI���G�h%Hw��Th��78�Ga>�W1�����N"=DY:b	�-)�T0zp���;��ΡV����W[QΣ�>V���,��q�Y9с�g)nSG[jL������yi��?ı���oL�O����78�MŘ��g��-cC
�v�뤅�oc��JW1"�L&mz[©>xA�礨ȇBjN����"���"ʃg�F6.|���9f4�\�ir���KTL���y���u�Èp|�.�& (��M��qp��3��Q�[�qG�k��j<�̮2��@A���$8���u��#1�"k� ��+6Fg��j���,���G{n%�d����R�"�NG4-}Ě ��p��7	�kju�(l��qCג��{�1@?S�Ow�F+�7+&�@U�:�D�.x��@�Mkʴ&�_u���L��=�x�B��p��3&-�q���0��SچO"��_Z�F���8��G?���gER�g�(-�V��IQtN�u�IH"y��tE�XƦ�7�us?��jU�>����H6bĵJ"CEh��c�M�T"��X�*�&�itW	��5}OJ�X=�08���^� ����q/Tx_+ZA�Cx�6aK.	�{����T*�%�y
�R
�@)��+w㺅5ha�u69��R���_��\���1��;\L�6�N���^8誏��(6n�j�dT� ����J��o������ H�`�v��-}7�"��q�|趴 3&���j>�e��
5w��0GXYΰA�J�i��N���oy�%�h~	`^���\�")߮i-J6c��a��.�}5�0���K���i������Ɠ��O��&��#�ۆ�\	��@�9�eg���P������R�@t��U �2� 3ɦ�U���,��(�϶W����1ar��!�_��D�xE��4�t .����a���=͖������W��Ls8������<��U�܋���q[�]te���cvA_1
Z`�]�C��xv��>����0��,��\^bf��������E����y�G#�{]e��'f�ȋ,��?l	C/�5S˞�&��_����7�/�U_D�8��~��y'��I��r=IlD~|���W��!����s��V^\�>��`b,��`��!]Hi�d���&�".��o�փ����x���_ߣJi[��7�*�B��=�������[��&pZ����Z8	�a�,6dH����~@��@6��E�7(H��g-Z"Cԅ3&�Ns75 D��&��}�� 8�?���c	E_3��[�6]����8�c�5-$O(�.L�}�tB�{Jӝx&$B#�@���T"�q�������t�A�+Oǥ!���dd@��\{&����Ő�b��<��G8��&]����H9#b�G���|:���ej�ҫ+��T�n�x�������*nM�����_�����[3��P\ʴ�E��;���p-�����
����A��;1��u%y?ʘ�JA�3A�!6��VM�xLGN���C�S)��a�w1�|�/2Z�!���.t"'�i�b����6才�	��,p��VC��[No���I��~�mMüJ�Ϡ�%�oD����ǆX�����I'�)8�~_�4b���%���찀�N��P�}�키��{����"u��O+���W���&:�,��,=}�������v9!�����M�%p��Y�O~�`����Ͽ�����.}��?��lm��߹���6�s(3��-V�#�U�\!k�aF��!yD���7�W 6>����̈���S����m�DQ�n�-c���Tf��%��ҭ��YW8*�#�wR$�,@| �*=^*{��;�V���H_��l��̍�2�(����9�<��kٴC�y`�=�"k�Ԭ�!���`sj�-�=�f�����Y�=�n�x���6�"&FW�z�gx�̆8�8�B��-�B�_��ňo�.i��f���?;����A�(��VԛqK�߫�GSx>f���%�F�c��Ń�A��h5�8uN2��}x�p)������j����o���Ԓ̳M�bY�>�᭝P-���d�B1%�c�H��@�9^F��#������<�8()p��ϟ����:�"���T 2<��ta�4�Vw����X�R�Q����J�Ћ��Ȏ��F�n�������+�Im��5x��ӟÍ�#��7y�3-������K_����~�ہ"l�^����n��|�k|b��A��'����'0s	���N.Y��c�0����՝CmďMJb<܋#8*�:��3�e�mi.�]