XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�����BV��m���X*��5��+��c/(^�@�}�U�� ��Q��Wc:J�q
 Vi}�7��9�X�tA�b;����4wJև��a��I��bRK�p���v6y�u�{���3�x�و�Ս J K�4{t�{����-�3&	HK�P�x	u^9�2���'���P9`K�'�胡I��vUK�)�^���z�����,�:�+��-��/q��a�E�$��rjB2 a+��щ�4 �p�!o+�@����� U26���*Y��?����*����F�m��~J��IM�7x۩,��[u6�M�IBFx<) �&H�t�Lf�IF���f\��'��h���+��4e�#J��Vod\�	v��(����`���#��l��k�w�񢽵5�8��7�]]�P8�Li@�P��"h�d�|O�]u��S$�$�G��K�`��qyҢ&0μ�n�r����;�VX����ЂFܤ<5�\=5f��S��,�wXG���F��v)�(HǇ��g�.�u0���y�<B���7_��O+��T)Rܩv��D���zM�44�����'ѐ�e�~$Ι$n	����"�;��^M��RБ}��>g+szڇ������^�f�(#�x;������=X������+F4g�`�����$�䒍��ѵ۝�fPhG!���|�0ᤄ,V�����X��_�J�$�����֏pY0�����I.z!޴�&���#����2�y���r3�f*�����XlxVHYEB    1377     7b0J�?bU�M<�'`4�}���蜥�����g�/C�F �]�rhäF��r���w�5�]�8�u�e���p��2"���D'J0���^����5��j���YL�!�?��,N!�:�n��g��eҕ��׀[끟��8ٗ��Tji�$f7���s{��J�����Dj�$Ol	U�]Ū�OWE3l���]���.�a���_+!���!cP������V(��&J��%��=�
>(�T����訬����|��}�@oy>�8�F��Q�3�֞*�	�� 7�m|�g!�v�U'`���j���ξ����,�U�Q�׽�Eq� /��OQcs$-ǖ�QE-b;B�-P���Ͳ���Í���ڍ���F�
ڑk�9��C��wz��¹�,�\��on�߀4y�y��0�+q��-K{P�C���/mY�5<(�@���Vӷz����5��/�8:����/4�X����ʇ�	)��א�9`�3W'��$��j�>��/nQ�{�_nzzғ��9g�����=�5A������b�8�*H��k�2y5��K�5g1�G�8�Ru�Ԇ&A�	�E� S�E�6�߽L����@����F�l��p��V��D �5ܥ���V�
�s�!�{�#�_`1˂s�x��%L*��5�o��$W^�d�Ƌ�ɳ�t�g���^Q'h��Ho(��M�����3�P���U�\>	K����q���q�.;`Վy�P�X�^�D�~}:�򓮟�C��6+�Ig��ФrH-fU��@�bD�Ɯ��y �b�}xDy�6�����"� �*]�pQ+�-�Q�zނ��bX:�����c,|#�'?�i�Q��ʲO�$rK ~N!Ο �H�"�܉!�	ԅ2���cc(�h'�Yfӓ��߂
J��Z*/����z��AQΨ���Jx�hMA�z�>���2gVa1<x�|(�߾u���u��Q3��=M�x�4����;A/����o�{�~d�؏D�_*���iȝ���MXh�(�Rqҕ�#ϋ�n���"���Wv$����[9�&,�%�9Ù������G)�]��������;�MVWX�vA��T�N2�0j\�C�L��9q]|�����@��+:9�}7=���z�Pf�����s�a��2�� <��݄��a�Tƃ7D�f���L��2#�鄊?6�࢛׀Uf��fی=�'ڑ {&�\�2�1dOh�B}������A9��]P��`v�l�;���¢X�b��$� �I�2ʻM>�6�������8�rj҈*N<hA��^���9 oLoS���H��Hs�7���ȏ�t)[2����%Fl�>�V+LA���pҶ�w9a89�r�B��˺�}.e�����5?g[��d��x}��	VgOU�m�y>�Z�/�u6�O����zM@yY�M�?����J_3���w�IC�<2�Q$�t�7���kz����\ ٴ~�2z��%��ێ+�
�&ޙ$:x�O�T��'ja��M��u��>�Gh
��C~]n�X�O�pa�|�������M�������'�nwf��T�[_�i�lD&��*Hi:{!�t3�C������(��G��h����)ɑ)֦K��ܲ
�� \uHF^���&�6��G�keV�����o��P)��b�
��Xd	� >UwIB͊�'���u˔��h�$>��vW�F���W��t���;͆�xDx���L��������Ce�꓁
�SQ	���)��K�C��w��s��]h�/zϽ�
�Y��a�<��?��x˴8C���#J�%, ���>q�h'90��1^:�)�:8�:��3tۛ�H}x�����m�A琭��# �LB��|��ԭ���Č�W�=��Ǎ�ê���w�sb�S���,x��(�-c^�������`��Q}��J̡!��`�+��f�tFc=���Ⰿ