XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����V�C6u(\$߇�yݒ��:d�����mu��\�r��n��o�t!��?�0ۅ���r֥̢�o���s���(��y��
�EDJ��J�s�vfO*��e�Lsg�[�&�i�?{�WWm~��c����7Q����)�JI���#Q����+��c�3�Ł��-2ey����a;�\T�-��ȩG�ps�A5��&	�hvD�ln�l�{dh[T��� ��Ȑ��J,R��Q�]q�,�1��<ˈ��E��$�U����Iɖ:n�)K^#Z��K{�M�\�,�Rm7�m�W��v��G�y�!I�(�t�ֈM������M��y�WM1�)~+��7�.���ĶS7�J����<�{y@Ο�.^se�߯�%����[����٘�9�tMJ��b#�~����c��4y��ϿyБ�&3��N>S��5o������,��j�W�>"��9�c\�ǒ� j�Y�����m������������hң�/�J<ru]���B�^@����{��v���RIu�z��O����R�QĈ��j��eya)��.cZ\X�����$�N��h���K�K�8�Q�j�#����0o ť�	�N���p�1 �F�0���?m�;e�Lp��qPi�����|��=��,r��P�j��_��$�{�Ts��/�����%��(�.���J7O��Aq5���W�����3�[&Z��3��*`4iw=H+S&YW>�:
�,�t�����F��9�3XlxVHYEB    12ee     7f0	M"ܡ�$N�fGM��G�V"�v��%�DXoAw�f2J���bC)z��0/u���X����7g⡿`�aOPg(iLYYz��%�s󦲇4�M\+30�
�҉�;�*���T�օ3����x���|���G�c��=v�����u�F��,�+�<�[�H�K,ډM9b�j���Ĺu���yˬ�6��{���9g�/��CdN�LW�΄(���
 �ի�U�U��ٶ���:�u!���=s���>V'
�L\/ ]�K���[��2I�;2-�X��3����͏��J������'|��Y3��@�h-��֗�@�{���Y7�(��)D�	�o�����~ ��E~�j{]� z�];ѥ��O���e{�V�J��j��A���J�D���U�O:�p<����"���H��	���[�ٹ�ͻ7uʆ8�|V~���3���3�U��g�ϧ���8�j������k�}��ޥ��ױ�e����D �m���Og7V�y#N"�\��!K����\�~%NT#���y|I�֯v(����|��[d(��)���bff�"�����F�q��؈t�n��/j>'������m�"��zIE�%a�	y^00̹�q�Õ�G�N��M��)��D�h�m=)��}o����)���U��
�VZ�z�F�u���a*r��:�Y���iX�g���(�p�~'��ka2�>��gs
KJuLzoB���T�,��?@D�\�/���QQ�{8I�q�Y���%+
�E���MN�I��Z��{�wI�bb�0�݁k�x@W�p�@z�j�SGA~2r��1R
��n�"�e���ً����"s��S?+J�Z���}%�ݛ���I�n�`�����ve�w#�X�G��S^�9NB�oy �1%Z�%�Y��a�g�l��Zī���e�?����H}?B�O�����6ֻ���3O4ص��L�/�l%��ƨ��JLp1!�G��G"_�"v���"@u����zv�ωtc��0�Vw*elĀv0��n�?G�7�Wķ�	���1K/�cK���8h�Ohi:٠�JOS��]�^���\�oʁwd�4�)Q�2F �N���ɀ���W�S!�Rs���u��7%�ߠu��W����"Z�I9Z�u,qg�ۻ�ԘhigOe����۴��_9�����&�_͛��f	��y���1���Qo�����ͦ�����&�s�\�N���=�X��r3ȑV�Ԓę��'Ŋc]�x�pҗ�4h���i��r��HW���;����?]��كr	�ǝ��(f�)�&Vs��m��j���o��{ ��ѝ��Y����h����Z,xG�=x�`2��*�Ī�j@�ϹȾ������ 3B,�ࠤ{h�
����V�ʖ�+K�r��#k�6lC�)Cmy����7���� �%Nr����7cV>�h��u���H�8�ė+�ŀ�`Y����X{����i�E�#�a�O��w�@)y��o�!�D�.�u��x��8��|Xڍ�Ra�ߗ��/t�t��?>�G���z�jh	����s��x6��`���r����92�q����`��^t��̧6�ѡ4|듒��Z��v��������7�O��:aYd�,A�F�b{b�D��f�;Y_�S�0
�b?Q�@��l����,�Z�T��I����)`��ݏ��ɝ�����5�+����8�o0hAc9�mHYe���d�Z�оŻ�;��B���< ��4�
�%JG�em��/�(D��g�[N���^�%��aZ�zYk.d¦�$7�7qZ�\~v�y��Z��c�	�SG^�ӲTf���21y�-���[ظ�<u=�����o��i&&l�/&�d�.�׆���
����Y�}��֍�����i�ӫ�Ҵ�-6�v�	�g�ڻ<�K4;�+@CbA��1�:�Ѫ���cֆ����s���p����r�:�8��A�}���	�°��H�p