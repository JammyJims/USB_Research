XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`ky�Ǆ�b���(�Wi�%���$"/�E��U;N\���T>?�u���i�s���M;P���W�6��������(�LG�g/��W`�}�0ꧮѾ~�� ?EQέ�偉Pl� 9��m�XB�p����r�5^�pVr߀��� 3�ќC��L3;�|2]B��>N;�pI¹�~�K��z��X�M}
^���֔�ŇDb��R���F����� �ky�;\��_�ֳ�H�f4S��l��X/Wϐ��70ѹ0t�[I�% T3�SD=B���(q�T���x6ITl-Ȃ!��mJ����g��T�#/4���ˉ��P�������?ޓ���`P/��靷�����d!�ȟ���V�Իn���Q��p��Cv�/�	E��Kh�է"tD<�^�g>7-'���9Pz���gW���2��_��S�|��_�5����Ly�������S��^Z�\�K�����Ƙ�M`�$HMK�u</�CO��ߪ�e�.���B��_,^Cb���4����]
��c�MG�Z�\�� ~e����	��y=����dc�����@?��_������8!�8sQmM`�Z�4n�2��Î� b�Ͼ�6�h���	��
�q���H�4'�m��6+h�ݏ	���f�����g/��_�]�8rq���_pgB�Ө�j���6�IyD����:Y��e�;����!��
�c���ln-����U�	0�.�a�=��7�]ˍ��u�XlxVHYEB    2910     dd0+��J0���vw����U����d�KA04ymH��+��`�����J��ҺĆ�(�����6��Y�0Ϛ8@�7�M���lxpO�`E���x@����L�_4/�����-���⥋$D�_,�lr6l�@�l��О7B�XP�.�[{
�x�LhrmD��H����N�OU�
愶��s�(v�T�&3��;�B3�"Q�L�l�#'yn/� ����l�F�,��:���j.�}��a�
�R)���S�^�����ѧ*���a��W��I�0�.�}�ԁ�@�P�;5F`P�g$<��IЊV���[n���`��"K�2�A��huIE�5w]�x{J����k�y��&��o���m����E
���z.�$U3H]V�N��������!s`7 ���>K���Z�ә��"x0�-���E>��DQb^�WfЧ1�X��.�-�󮂲:F2�t�6���Ͻǵ㗸��"�����<gf9�E_gꪬ�Y'�]{�\AD��lT�������1S���hOm:��z�+����>{f� �uaL�8���+\�3%���(�oX�j��#���x3��J3y�W�N3�,�q񄍸��!X7�7d@�)y�1���9"l��U������(������)}5�Q����)�K�nޏ&Pn���	��f�\��f�ܸ��iN�f�!����ܧHT��.�b6�����J���V�&�{�n��O ��k5�L��i$q�HH�>b���F��4����K�@�$7K��F��T�¶9���?��J��\Ж�:	�8޳9�=��Gf_����50�vg�°�}OF{��U3�4�F�y�}QFB�nbs����o��IR`�����ć�h:<Y�4O�w�B
j?J,(r��� W��n��4��>��,�X�6{k�%� �Q����$��R��ʞ�s�`5��n�,l�X��H?�`���|��6(�ڗΓA��Z
S9��B��T�͚����E1^�+R�pY���O����^�j�ZC��kWU@�x�[�^�Y�d1�e��	aKg�j���lGI�nl&q��F��/��r����~�1�0�`(���=�[�]A��`�d���C�B���ۼ��bC��>=�К�'�����s~KgǌG�g�W e�8�qp�F������ۮo��K��2�o�� ҡ��o�ňk�,��d.�t��i�V6�)��_�vv�ȴ&��cg��k�@~`��Bs��C��Đ�[��3l�f��02�6V����
W��jX6�ܨ4��{=���X�HSд��N~i�
��z�®�I_�t����c0�5��,Q�R7y���ؿ_�R�o,�5b��M�)�v�� P��ל-W�|�}��rI!T<(�Ϲ����)�8k	8|Ȳ�%�(:Xƻ!V`�.u��Ul���CB�V����K���Y�Is�55�Qz�*���& 'no�,�&�쩽��n��������YL1-8���H�䐏g���ꟻq=g_'�H���!9�O����[5�q��-Āk�ʱg���|�V� ��M2�X���T#{>�x�ӯদ���v�&�0:��V
���B;53���ϊZ�V�t	zA���f�a$Yc='.��j�`A~h��8zQS��m\%��!~U%$,�B[.����7��eV9�#{Q
Q|l�Ʉ���v�V��{-GK���"�*X�k��@>�,<K�V�.6�~�^/�`�!��w���O���JN�Uɸ՝c�WZ�ʝ0o��&����#d�#� ��{8@˺n��j$9r��Cg�$ұf���X�\��}Ɲ�yIMA%�&�|�N�W3�҄E�ӑ�):򫦀���N˰�J_��y	���՚�����ّ�TM�g���E(��}Y%v��c��Kq�Q��xC^ͤv��R��t>��b�67��b��=���]�q�e �(�����C����f:!Y��6��c7]��hxچ�H�\Cb%NB�9�q�B9s���_��J��o���$f���<8W�@�x��.�@�he�0�.j0F�2��Y����m�g�tA=�9o�B%r}��Vu���D�n��q���Ƙ���_o�E��~�w����?�^�&�}Z_�z��Wɱm�<�[�9k���9�;zT���C	���ģ[�GLr>�[1�׬�;��' v��{@��&����\Z+TM�~��y�=EzM&g�E�<�|����'��M0�*��N��^����I �NvQ��u�K�i�����&EȒpW%�Ӕ�M6(i�<�/Pw�xV�~Q�u]�A#0l�?�-�Ʊj�'"���x{wQ��"C��!�D8K���2p�,RԣRH�Ct���*�؉�����̭ies�MEAB�~��e�L���Ft�?u6�_�;���c��4�/A��oo��G#yM��eD�;񜓈�2�c��CN�ەƗO7w�x�r8G���SB���%��'H�c/I�hxp3n�*ɤ��;9y�	���O�͗�����`�)`xH�J����k��Eg=���3^4�]s�$��^�ʥ�t���鸲f *�,�r+PE�%Z���:�R.��Y�!]F|� ��9��X��;uM�Z2��[�V[I�O¨ECg�b��&��-�j�/잩y�}g�������4��9�B��nD�Xh���ؤ��뙧�&g�lfq7K<b��7�:�	���IR����c��~�(��$ӌ�@s��(gT9�nO����U���7{�i*�JJ�eb��]=sr� Q$���9�c
EKƘ���y�W|Y�X\^��
/�58�T[Z}�V���6H����_º�?;�GX2��O�'�v����������!w����Ad��3a�!i\yG=;0gk���Lˆ��E�I�)�+��3z1�U^����L�
�<J���b��_zh�Gp�w�6Jo�����p��Ӱ���y�z��T����I���U�if���Ȇ�쏣��^�#i�0��J%Y Wޚ+��f�H���e)&8�c�	��Aш ��߈�o΄2g�#Y:���7�ql�j���P�ѵ���u0�<���n��7�\<	�p���{��]߮S��QI�b:u\bLVq�*�mA�
��RpnX���I8�����
ʰHK��#���K��v��Rw}N*gD��5#���b]5����r}8P@c����g����]F�./P� �r�4��fZ��KkLn�Z0��"�|itV�@v��O^^5����Bܩ�kwkrwF������V���v}}6��M[΋%~�s�V|蘿N\v��e���!�A7n_�z�������?����Wp \Mp��mf/ɰU�eǐ�LD*B��5���'�Q��		�iK�j1�z7;_V\\�N�g���_^�)���gر?ѻ��?�rk\���BR��ղ瀚o��pYq�F�F-�