XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k&@�����-��g$�i�U�a.���m���X��mwK\w��B�b�9\��  ��Kp�H.5)��_����a* s�̩��ʁMdRl<	�>R
��i&�/�OA}h��BT�-�C&�G>o�O�pQ���a��a'�+�~�Χ��.$L]��o�W�)J*Ɩ���Ռa�o	��<�X�_Q��@nQ0��)0[�O��T�+`�#Y�����I�x�c@�%��5��鴑�|n+�׎�	/���|��+7(X�0a2���������IR�{��g}���O�y~=+�ӗ�5/aU���a~׹;���s���2�cj�͹�2ҁ:+3
̪�W�|K'ND��g�N�)��>G�؅n,w �<axό�?�֎��u�7�8*���Ȁ>ݳ��0y�S=▢13BL��J�3����0�9�S������ D�ح�>�K�����@h'P�)Y{����/_ʺ�!&?���,\��}��	2��U�.��k����2/Z)��3B��1C��hdZ����ߟN������D!3Ő۞E�8?�k��>��#V&JJ��<p�́���&����_�bm�I���c��p9�>թ�i�0w����D�6avF}Z���~S%4���#a|�e��>�<.���(�V>�/'���0�a���x2ϒ�c�Т�7�����U�S}A�hG?\�*�qa����(	|&�Q�j�;f��9
	���m`����)^�l/�%-Au��+z�9�η�Z��V<�ĨB�XlxVHYEB    4395     a30
�W{츝��P2ɏXW���+�n�51���4��R)21��5�P�<��兔�u��C�̵���V�[M��������(v��R2���4C�%m7Q�6�H"�93�*6ӏ���f�;k��ZL��2�Vc���� �m�bd3'�B�}����~����������]2��K�~(��>�
�T���8��j��}�\��Ɏ�+_FGgT�xx��=�ō�?��T�P��tqm
�)4��'����]���V��2t���4�;Z09��s���C��wx@\Xr���@̱�E���J�'s�՛�=����=�K	8����*b��?��i�q�1���ưQ���
W7���L����aL��TmD?��f�F�g}� �A���#�]rֲ �[HbB�ÃH&p]C�b�D�G��IB�?�ZA@H��&8�K<s*y���@�a�j��;��X��� ��#�}I�FĞ�<��+H� ?�|��ܒ���2Y[]�&���M�%L��S^��f���u�Z��q��'���(�Ҹ ����9��
�<i�'a%� m2B�_h���|�CK�hH�%^����2��hq�Y8���<� Mg<mΈl�ͯ��Ն��jBQv�7<@|�4�)Y��ޘ��+����\B�3k��ݓ��/����)�,��h+��ld`[f%d!�cAR=ߊ��&k��d�iv��!�m7�Ѐ����q���X�Q+K�ܽ�"b(�nH�.�:Sdj��GZK&r8:�W�X�Id��W�ҿ~���u�w`��n�y���처�7$P@sC�����{\8D<=�>�|ʐ��	z
5[��Ѕ�5���n��(���xm�;�V���6HZO}A΍c���P�j²Kw�;v]Lꟙ��ھ W�4�6����.a���Ila�[�~�$��h��v�:^�(�p�'�g��`mMh��j�*�c]�T��Օ�I��H�`0������"O��5������s���=,S�Q;�4�QY;���P��4p���L�k�Cа��,tQ��%RJD^���0(���}O��-��{�k�����oP���;��� �x����=�<���0T��V;>�R�HZM��_G��s6�X��ŏ���A�� �hr��4YO�6����Ԛ�k�&"��
��G2�dµ�`�O$�_σ����<ȍF0Lb�	���Ű�����)����E^G��V܆����o`%��Q�����U���m�hOe�Ro6�N��eȏs���\,������XE������k�[�m�*�n�����B	����k����3 ˮ��@]xgZL�M���k������]�I9@��8�\�?��n�=nm��Y6�P�����k�٢ħc�� ��"V���sWvż����|��,8=߁d�6�sv��3O9d�$��o�����&y��1G̶���BO|�Q��k42
f_t�/�N��J�DQV��ߨ�?�W�� ą`^��OV$�D<n��D�'���מ��;�D�;��a{�<�Bk�ª�M5U�ƛ���`�>��-:��~g��`��ڵ?,N�4���]4���椐��dN}q�CG&�wn�ĺ4l�}��(.��d�3G�KMs���冹0F�M�=��M6��Y4uy�^
�Ɵ	"M�J��Fvvrǭt����$�������X��Q(�߉�>�f�(�`C�>�Ԡ ��k}��pg�mj��r��@2H\�͑%�=d���o��%��nC �����O p�1�ޯ�ĵɒ���_>�b��",�J/����Ո9�a��Q����ċ�B�VF�N��{�l3㙙fAP&�x�[T�H/��d�e���ᩙ`��1���G��IU%�E���N�q�_₽t���� �"�䤗�5W#<HB�(l��oy=����/�``86Tֻ��nLf���Ą��˯�8M{^���H��b-�&ҲU�p����3Y-���V�Գq�]'JN�9����7�O��8�M�	
]7��#_2�U�v��/��(~b~zE }s0�ž�E��F�����L֤�ý�XԞ���1V�+5nUP��v���j����w©	)6$�bQ�E����	H��n L�Z��\��/T�u�\�]��dm���-�,t� 8�&��b9����{~.ȸ������o%xJ�Y�Z{�1�=��|oaWS��gcg֠{�h���ds�/�\5<�Gr3�k1�X*⮼���~��O|LW���;�����5b �0h��(rͭ(4�~E������k��m�7*���#��˴b�T64+��C�u+��D�.	
�B�s��n��8��8��f��-&y%Ā�S�ꂼ_&�����`������fm΃nfP��V�b�$Rׁ�Kl�-K�v����m�YH.��Ow�&�I���PS'���6l��a`��'5�ˉR�����p�~(�ԇR��S�����TV]�������`�@��ףݝ�$܋��#R����X��Ȕw�$���<����