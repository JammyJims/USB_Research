XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����(zfu&�� .s�>�����a��a�<��O�:sG�Un������!@�3}�΂JF-��V�+d�=�_H#�ev������/~h	\��G��IקJS�H�屰�31E�?K����X�VM���D!��� �ȹ�$$J�t��p 8�,ѹ~�@,j�w>7s�&�e;�c���('P������ {*\Y~(2+D�ܔ2d*Y��R����>�d�1�{U'�	g�f�n
���6�?�ѡ���kS�{at�da�o`h	���Ѷ[=&3������1���D�IJ�|�GS��ZuP�V"ID٫�g�p0�{��#�D��	�l%@��ƺ�S�ڇ�ȸ��z+֥���$����0�{Q�(�Ǐf��B��/��^?րm5� *oBx��!��x5��,�6� sDe�����!$t׺����]����@ؘ9������)�1G�R�9 n"�s��50A ��٫�9����􏏮�:l�.�	%��<4`_Ö7�enO��)��/0�~�!=��RS�سR�x*F�� ���|�^"<X�+�����b��h������x��Z���J�GC[�~1c���ۃ���E��=���z�W:7a���H�c� �8ui����x �Mk��E��w��y�H��u��ΝҸF��m&|�|m�T��D���'>��w���4�8��zvZ2�)I4$���!pl�J��ơ������"�O2�6��1��զRρqc����XlxVHYEB    16ac     910-ّ+�e�f+�#żD�k7s���`��:��S�tC{�䕳���=znI�1?�D| H�� ])q�X%�e�5���L"���ܺ4`勯m9EA�ɧ',`vr��@�m�L6;"5��̌Դo��	�%�9f1�b��.WL��'㎴9�:6������`c��Z̥�9��LA���Vs�(�]�w+#M�`7:FiC}f��0���ɞ���������,�R4�W�]Y��e�z�83,���S�v+���
>��cѤ�U�X�}�=%-�I�E��V�I�O]]�!�a��n��5g8���ւ�b�+ř�G?��t&6�adwx�4^��=�64�=���1#�ߌ*ҁБ�R�}�F�F�8ѕ���{�l�Q���
l�Ͽx�5ID���6�q�#�eJ���&=���a��(>���%�>l%ӹ��U����::�"����߻�A8Î^�%�M:�)�޾`	�K�l8�!�.����WBq��]b����=�M�`�bA�͓ڪ�*5+y��-A�kT�.�����^)�W���	�zPĀ�#3�u&��|�{)z�O>��3P�{�olx�G���$�kqP
6��m� 9���\�ɤU�s�:T�N�oWdK[[^�#��?���Ez�����dy�#^�����ڒ_�3��cG��y�6����]�߄O|d!Q_
������7�p����ⷠ����&�#_�tBϿ�dis��)$ᖶ�١L�9�ۅ�Z!�k�`O?�[��F�>����?��b�X�m���v�}$n+l/��=8�	�	���؛C��2g���qB:���]A�^��'�c(ΈjX^;��������E�Pbc�Q��>k6���^~�"��o�{���`y�"x3L����O�V�^�nC=�Re�$տ�M����)�Q�0]�'�Ԅ\e�1�=r{	]�+���;��Yc��U�l�T,��r�F�ڊ�>=�f�ds�Q��c��}r}4և���/��]���5I(��۬�	[��BɁZ��_5{.�''�R�/����Ai`��@Q77Y���M���B|�|,����?���q����GP@1Y`f��Ϊa^�(���WyYUXq��o�2{�n�7B��(nt�fQNV#�,6�`�.�Hd�+�fI~���"U�������k��9�y
�{��e~�Bf�b\��ޟ3!%���2���Iٻ����0�y�[��
��Zi%Ptͷ��@щ��ܱi�D���W�F;�t�I��c/,=bg�{@M

��d�G�R��B᳞��pH�,�������@qE����Srg7zrC�*�$��ݦ��-�/���@����Śy��p�L�j�joR(ШPo�ѫر��7*�3RR� )��p\��+����pN��3���k���&���ټ�j�u�����ï*�]0Z���.t��}$�t�M��^�����B/.l�7���Ӓ2��4v�{G:��{T骇ܹ'FzN���U�{�K�_h1ۻ�DO@��B+b�և2���b�[�ٷ��T@���W��7{�O��������?���kxkN,�=L$�����9fl7�iѭk�2H���[dr[��[�CR�bY�����
��u�?�h(��̳gΕr]�N(��P� QH���̹zrZc*�kݥ�pk2���3Cs�Sw�tM2��/�U4�B��Wf�w�@���a�D�ro�a��1/h<i\���ޥ����ހ�)�%	D��{a-��+���>�nea���
tT������n�G�2���N�������I�+Ƿ�N+�VH���FjR���	�M$��)���Ιa�5n�p��HA
<�}��=N� a	F��B@*��Ar�6H`L��?�aVu��� i>?Q��Q�Q��ųF�S[�L��;�	�0��h���-r^1�e��#M�/�a8�,gll���%q#-{q��I.F���h/�N�����1V�2�hP�¢�'Y؉ۤ_��=g�p��=��!m?}�	���O�\���9Ԫ���:l�5Sl��x���'���/���42�~T�5��,R�' U�;^P��s��Z�*%n�|_���n���"�9��>v�z��4(E��g�D�p��/[���$؂k����Ә�Y_=� �I=�%���F䊙�e���~�m��x��,��ejs�T����t�rt�� -����nÔ�
9�Ǹ-1J/j��nuP)� ���X�ë��wߺ^R|���HlI
6@{���䳙�X����H