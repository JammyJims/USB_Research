XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k	 4D�E�|P!�|�*Ƹ�u�#���d�R�ik�O����|�8�i)7�9+΍��d�Q%�-`t��qȖA*f�{�D��A�$|
ưF7���?5��:�/K�fK�0�~植mY���6���X@bu�����W9��	,�����~�M�ŀ���O�!sK�*��ϛd�{�ʛ���"��~Z-bJ"M�  �
蛉��3гUZY�f�u��f{}��ՐJ4�!o@6�!��Uu
�PZ��Ay�D}9wq�#�%:�&�Μ���:�h�ɧ���%�]�裐�I�p8BkM2����,�w�������Hc�r��7�d����y3�`��6HbT��n�t��牁i;x��	\�^�nY\�W;�w.#���נּ��І{�n$ʃ6̃��պ+$d������k>i/I4қo�M'<��pW����!�����hǭ;Y��{����1�=�[s�����̀�[��� ��=0�[�C�:�p[ ?>m
U
�Â��C�8�Ļ}�mQ�"[@�S��5�Ƥ,��S�������g(����ۚڃ|�6J�.�_81��	鿉J.�������q{�."����₋o�k����).y@�c��7S����7>�l?���FcG+M��}X,@�o⇸EC��u�Ɨ��*$�'��ڑ��F��I^��z*�~Fܖ��a�W/�_�����V[��!���$|�5�@v6���Wx�;���Z�J�"__Z�F�
�{�y[>.�a�X" !�i��dXlxVHYEB    3654     c40?m9-�kw�|�1�v�O�h�gH&��z�@0W�{t�ª/�g����m���<R|+f���z���qil��p��>#�bo��\���g�.�	�}EjY9���V���,�t(��W^�_)(��M1��?$͌8`���s//�ԒfW��@�ǣ]�C�PR5��γ����b��V�c����Wj^�x��H��G|O�M�;�W�"?'f��׷���
�-�+���Z�Z�>l��'�̳���%2���H�?Q��+��)�����/yٮ4+��Z���J
!�gB�g��hF�'����w�π$z�������>fOt�R�J�4���Mk���6Z�E��^8mD��/���5V��;�������SK=�~�G�`d���>�F �g���3���o�AyiM���h/긧
^���o�}�w߉V{��VH5�u��go^Z���N��4�ؠ����o\H�[K�; :��f���M�e��4�P��53%�&�^�ٜ��`�a�ek�˛�E��墟fB9��٪<K���zb��˕�H� �i&��(��͚3��s AuzE��(�cC�c%��ݙ7�R�\��*(�x~�:���^���3���>i����cm��=�)�IT�d�Tu��]l�Zй+X�B�|T�YC�����M̭���1�<?���G|��JKſ҄�/�F��Q 
p�*�U�mڲ��)j�n�veI"/5���s3P�u�vhŗ`9����0 �ciU��x�5C[J�f'�D��9��R�WEg�Yf9��Ɨ��1Ry��fT0՟Q����f ���c"�E������v��ċ�N��[
����L�[��=���7���g �d��x�45@��-��5y�n�/.��l�!0П�I�� g<�a�ߛAoX���M��@°��6�����1�*|��!�f+�_Ѓt�9�YJv�]��:����p:%��<����H����cň{$����޳YT�|�;��;�ٲ��I�EkՉ����W�8ϥ�!k
2ߊ���qUt=��vd7q�iD�d�1])1z�#��)?�FȘd�L��n������\7���,-t1�,� ��ӵ6�@`�=��q.�L�����r4����u����1�����`%p\(�}��1�͂��2�8�:]r]�fB�KTt�O��櫱6%@���u�9V!u*��g�Gݺ.���݇�c_@�	�T^T�+�f'&��;K���sN`��4����
��mM=$K��w�wim�2�vŻ��"��
�NQr�bn�?<�C�� �"x�έ�9Q�	���KN+��p����#�*�+�7�mM��!E�6Gt�?��P� ���k�Mc�`o�J_D����zŌ�;�(�Yo�cW|�kk�
xs		!���y(�:���h�^�����eJU�!J YJ���Z��	��`8��f��T����K@���7x[7��W��C ��Ͳ=HƋ��E�ma����.��	��$xЎ���16��QѪEߏ�!^��{�-�U�0�/h��
�������0�Z���su����������3���!F��u��kwΆ.���@���|֒��d%x��ۮ��C�&��: ?���E�ť�%�ʖ�w������ �Gw�(��A�T�9�Q�hC �J�����?�h5��KK2�ky��ݶ�CD2��٥t&Iɒ-�ŵ�N�e��s�)8�{��������Gj �L|�P#I���T�&�>,\�UEZ���2�D*�"���y��"Q(�w��eT���v�u�A�]	r0�f�R��]��ɰ�$�B~m�_P��Z?����Ɨ��Vnok�d�����^�P�I/�s����bZ�?U[	���4�@���#��g�t�wR��R��T����)�\!��dYr������z��*��D0�A^�<,^]�j��&���<Q��&A�[`~�����mYv9�+����.�u���0��=�F���)ς������m�n w+��NHc�p�m��Z08�3��q�2��5���t=�Pc�$�s!�AW����
jo��-TI-�M
�Rʫ}Duz�7ݘ�R��i �d����o���kl�1�|�P����Ը�/����G���gw����t�愒�iVi��Q�T�o$C�S"���+�zA��0�� آ���A��
!}r��g[m)2���b�����%����*D[(LĬ�%�Mn³���	������.ɔ ��q��?�dd"���hPq�.5p���_N(��Aj�:��䵟8zQD�En��4Q�-v��΃��L�ۤ�;�����%�� �t&�d�F=�W%7·񄨛ݿrR^��^���/ �n�(��"9�3e��R���D����i��8��t����L���=�r���[|w6�8�E�/����$���ڢ$z���^Ѽ�B,�:�XZN��#׿D�T.�/c�ARK'����NIe�f��P��8�TB��>�x"s���5��|bI
��/�P�t������-�b~���<0f~�֫qr�x[_�%��n���qQq������-��(���y��E�@��S���e���[����%��Y,����K�2��d�D�V�q�-0���e�-f������ǬbE��5��%<F
t z�+gM�3�����g(����в���Yfų����ㄴݔ�l�%5���V��w&�}u��fd�6��3-5�����s�HGсc�����ڤJ>�O/��*��Ox�-�1�`v[3������hY*�v��,o����O�W�0�E5�k��,�T����r�LR�u�� ��,z�,�m�<!�p��aM!��4-gt������D�����t(��'z����`�˓�x:�?�ogD���i	(<$�M�t`%�����|Nɥ�#1�^���Q,?�Yk.��
�>^�JH��m;��rA�����	�}
M�bb�dz�T�#{PU��+N^���L�
��nP�0V;l�=�~d�)������d@7��8�t��9Ђ_-��<&�tXOE8���Ym�@=�\b�<\�WI� ��i%~�u�W���&��T�[�	��p��