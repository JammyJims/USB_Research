XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C,��@��<8�'=�j)/(=^�vll��oZx5]���Zr����}����*/F�,��N/����k��y�W?Z�כ\�5Y%��}P�H�E{�.����IJ���&���
����3v�U�+�w�z"��g󉟸�+U�M�ïW����T3+w~�����]bξ��ЩC�U��Q�9�Y6�q'������+ lپ��d���m�ᇠ*�&��N�nG�7�]}�x�������Q?xf\+mrc�g�!@�N�A{��4y�8��5�vZ�����$^��ɲ�}@�!� �F�9��J�EB�Wp���2N��ݟ��3���֗�5}#�͉Т��ږ�)����'F\���ԹLH��h�Jp�~8d� 
��A�vG�.��U��dG:M�S|��~Z�]����ٷ$8��9�vn��;� 	�CD�T6Ud�*�4�I*Y8ȷ�Ų�&$��'ŗ(��ĸ�)l\�x �BgYg���O��(�!-?\Ihfm�k>�Y ��N��]������)ܖ  �5?�=�p�����/�� Dt95�b/����ܼ���4�AT�$E�X/"��'���?���1^�L�7m!�Qv���-�4ِ�"�z���qw@��4�.���_�V.��,�,�+�at�'Q��"�Dg�,M:���ꔳ�@��ktc�N��ib��諨��Y��B�>gW�����@۾F�o��̀KL���4�����*Q ��s�a#�.HCi���|T�Ud�\:�7|�+sE�4�	!�A�o���XlxVHYEB    2b87     da0Px6��\#�&�4��8Q9���SF~U�3'�b�N���
9H�|��ٷ֍�͕�;�y)�zk��Ȇ��q��?��{@�
�Y��Z��}?�ga�%�m��<������Y���+RY��	�Aη⁋2D4�-j�.d�+��L}�ݽ���.��mh1]�d��O�P�[;ΡZ'bB,�l:�2�\���[���/�iJs�Lx�*��͋'��=�� :'CgF��I��E��浄�l h�ڽ�i�ؠvy[m�\�?핵�ؠq*� �銼��kG@�|�2X^l���*�b�M!?6R7�P��<S�Z�����V��B��5z��������������y�̄9����'��A7�����zw����>P��D�G�3�W�A6Y��~���eM���JZ��3��9_��K�}��K�8���}�y�Z��u4
�c�
^4�h"TX�a/�a�9�z�z_C7A��dkώOn5��M��g6�M�v�>�q �:�얩y��H.:eo(v2�/���5��i�g\�bj}�WqQ����
����k�3�l�t�x���Hx�f*��NǓ���9B-�JYo5��!��0����q���)����ų��W���P{��U���R<�w��z%ܽ�c��L}��l��U��9��-��eP�����53�v���� �>W<Ӷ�}3Z4��d��@�-:�!�
�i����|I�5'PDvb��و�3U�cс�bq"dR�����a���}{��ewQ�o7� ���;�d+�I� q�̼�8�7�N8#� R�J��l#,�ҧц�ۂ@rIOԬ������\��w�K"'��~-�EvqT�8��MD�DGᷲ��3q�[%��Uz�kr�=$� �)�%'U��]��ǘ����Yɹ{i���~2.4�``5�0rx�2 y9Qy��ѿ�*?)鮟�?̻̘c���QP�^6\a���Tl�M�ϔǇ`�GI��%Ȫ[L*j�*��o�����	�]&`ſ�y��TaΪE�4��?���2����^ �xt/�F=�u�}���6�\[�?\k�o�܎Iו�,��=�6�&�
K?Aq�=C��Y����ZD�Z�z���#�R��! �m� e�<��z�=�<fiҥ��>t�f{p��Up�J�A����xª�7�=`����)�T߭�̙7��}���>�����#�w���k�pi5=�	±�o�Y�<�?�
�����mA�
�/=���H��	�(�U�\��Cp'���9[�if��3�]��$���P5�G���-VǪ8F��O��	��8���x�k�7�������MgC�/k��¦N�p��7�-�����}����D���Ą��$������?<�vK\"Oܸ:����Є+4)�((�|�B0 ��@GK[�)����e�����<�T9�É��y�a�y۴�5=o�%���W�0+�%�AE\om5��M�w�$�j�ڑZ�m�[oEW�u�E�L{i,y���yּ���1�Sr���2��ĥs�ڲ|������,�#���z7W�~M��.����'s�GTD��놛�g��W&'�&@�e��ܞ��t��hrQ��}i&�/		�F��y������^�O�,-�z9Q��<�����MT�d���>σ���hO�-�����b7��ݴ�˵�5���Xa��������!���4���%`���+�d�_P���ajO�,A�XZbqA9с�=	�I8��/ޥA3���T�7�M�L�<G˯9&�{����BD�9A�"ڰ���[�;��Q��ez)��x�x70o�K��� �����dN!T}z&��YF������K9l�^!��Ӊ�^��ʮ��Z�nE�6���(�9�sXb��������u�"�P�t��vY�8f���+���Tu���p~ˆ�,c;X�zk�6�cI�i�]�5��� �I��A��(u�f�R�WA��	l��)V2�a 0�/�M����:sl�N�27γO����3vȟ��Fp�o>:�U���Ǭչ����oo�F2o�{���k-Tڣ5�W�N������jr&P��^�tk1>e+�ư|0.�1ˣ���I2��kG� ���K��6��d8�F�N��8�p�9��3�+�{�|�`p���<�
�a�`V���sV���j��{js��g�]��>T}��PXg��1��P�	w�X�E��<2���蒡� !��?J(F���'Nw5��K��
�������0���Zw�D�@�=��(c^`G��B�$��I��3UMPsA/k�̂	R��_wJ�
�}��'H��10�C�g����U�6�����:Po��!O��%���:]-ģ"|7�3�К��\���<�B�?6�Gs1C'0-��[�-��4){翖�7�F0��0%��4d�?�x�\�	��ҙ����02��p�k0�z`8�ϛ8�7�vCv#&23Fkz\��P-�<v��l�x��r����V���n��+� Ň3�[��0�N�_L=���Oun1 YM+n�Q����qER䱶=�a}�\X?��J=�w*Hb��s(����gC>���N:~�x�|a{�f/�8,�e�xd�a�тl���P3�a�I��^5 ��.oM��޷�W�,Y0=����[�Ж[B0H2��vD�����~�5ד<�m�x�������F�g��Dʏ�8�*KD�D/������k��������$Ɂi��#h���p-3��������X|0�?)����P��t����$6���k2����z�5@�X&>�������n9�/���e+��T��t�28���}��^x�U�h42/D7�Y %m�y �`X�fĭ��R	�,�ER~_}�%/�!�H�:�a�ڥV�ְ夕g%�z�x���.�ba8ZJ�$�.��C`���2Ѳ�_+��h�'֛$[¶+\�[ZL.�pfа�0�� i�ެz��:b�I�\HiS� G�r{��z�Έ$��9��W��K��6`�����ű�x0#�Y�i� >�e4"�
��&�
�x�ݼYi��*[���9t,��_���ٽ�D69���t+�ý���������&d���	��A n@K�9[�>����%��el��nd��K(�&�Gj}��OZ��"��a�V�Nh�d���W�5��dO�� �O=�Rh���g Y�'���d^�����9`��~�hM�5s��Qa�3m�M���Ɉ����Zk7�����G¾�S �1ʐ��%(�����o�.�
��7ү���"�M'�f� �7��:�'�)��H�L>����Z,�0���`;�'ǜG87�Z��-����VLiP��jfo��<�������g�>/L�tmS�K9�=׾Φ~��Cd�W���b���s貈�:��?�ň�