XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ؔ�����|	���6o��΀Wѳ_�0L�;�N`� ԭY����N�o�Y ��y�PE���B�|l�j�����'�HzF��f�����]LȺ̡������=��nr�H�zW�0oې
I?UЗ�75E���.���đ��$ ��:J/G� ��x�@����G������(L����\@E�a%/�BOS��-�\�))3�3��3W���8�籓l�pݕIv�����'`2�k�x�X�`��
�^ۇ��F/�	��!K�d�_�x�%~�!ӏn#2����B�)ҙR28`����=�% �Φ�T��=�Q8��o���,ґBCw�H�Rɥmq �%��9Z�T�;�P7�s-|c*�bw׷�f������b����<�o(�S$�j(*�� ���w�/���e�>n��y� w���-�G���Haj&ڏ�r���ղ�u}%�OSk1G�dP5����>�5��Q�Ϣ�]7�0�KŁ�1t�'R�����4� ���"-Jwm�Q�}�#1T��:A�&�_�3+(�H����2ӷ"�u3���'>%�P��I�?�t���1X3�2G�+����*�D�)�����/��%��;�i-A,Ź"�kj=	a]u�k�Ft��j�XOӏ�T���h�E^TX�g�vĬ+�e9��Ɩ�?�I���)�k�?�����~ۈ�џ�B��+�՗�s�諈��x�l�����G����y�f[�A�ÈAiobR|�9���.���(��`��XlxVHYEB    19ec     9d0���ޫ@�n�@��}�K����+�Cӏ�]�����M\�$��OX�tS>�r���M�]X�>W�ld�M̢c�jGj�v�It� <��/w����'+���8�8�d~Gg���5́�O-˕�xi�	N���W�W�n�ʚ�@7�F!�sհK�}oJ��z�"���m��Rߜ���f!�r�N̿�����$)�k�B����:#+z�F��>�96*3��!��|�Dtz����F^v�$��Z���8Q��Դ���H��?�R�.@R�}M���gώn���hn!��Fއ�,�}<��$��1"(4_��9̷Ȕ���n��v
���Y��4Z����ٮ&	B�0U�F<I.c��f�)�Վ׻�L���GM��j� ��&��=n�ҫ?Ļ���D�y꓊L�=�� ���_�O�C\c�<�hT�&'�WYW`Ꮫ4@@3�qs�*�>�Q>e}4��L�ip�3δ����0�l)S:�X��"y�j9Fj���Dl_�X+����R�wW���P�����o��;N)�t�sW��P�0��=�d������bXncGw�!����K��|V���3k���F�+&���G�u�f� ���^j�u�bij_�Q'(��	�aG:k0Ɩ���jUʈ���I��mRs2��9��Hp�Vf�&ٗQ��%@��~:�O�����ڧ��'���I����(]|����Q�-'q-����\����H '�Qb�y�Ф،c�b�Y5���M�Z;ꄻ��Y���/��o��m��Q��K�Ԉ�8����𼀑Z�;�>�ZK�SgEe�F�cd�?��H�a����!�JâN�F=���I�k��vOq �o�Ö�9t��b��Q3��g�n���rPJ�/2^�i��N����b^���q,�4�87�B�]��t/d��_m\�	��Rl��(+�F���-�����$Ғ���H8�Zf��\~��H,�dvM�f�HB�*|��`��gc�Ԃ�*	����t�-�5��/��;�9��iT��
��<F��Sɬ0<�	�z�a�v������6C���f��1���ۉL̲E�T�x�o�̹��yC[4�fU���=��	v�R�3��]�z�n������(�}���i�U ��b����I�<g��'�����3���0k\Ȍ�,;����Q�H�7
����F��T���3�)v	�w:ێ��ʴ�u�)~��(���$��.��q�Q�/c�~d�Zo���.���]�п�h+g_(��!���q_pb��[�&���V?8υ{��&�w�,+�B7���?��@
>������3|��a�N��_���eٝ��6�<+#I��=47e^�9y���� O���O��舚�c^�GnRW���_�a%ev\���Mֵ�n�������C��܉���K������=���R���v��� �D��,���*T����Als0����������}~��\Z(Tf�K�F����C֧�f^����U�~d����k��|�A��M��!��ٳ�����Ak���NfT�l���2����H�t6]/�;��0���L��@���g�bRURC.�2ƴ���h�,���E�H�Ĭ��v��H;5!v��j<�M�������+����3��+1,$�����s�2����q�8SBo�0���^۸�������C1Kh�$.Ox����杞� �g�{�����t8FC_9a�|���-�6>A"�r�O9;��[�s���g�L��ŚV���q�Bi�+j�8y�^� }�^(o�9�;1��c,!-���xzTq��O����`O���P�I>�������1*����(�1�n.�WZ��m]��{A��공�k��$b� �M˟1���k�y��M�S�:{��!x��
n͘��k����h� ~Jn8�+l �8ϟ�݂��[L�76��v����4�$@��< ����u5,�X�ҹ����q�P??m	�q��	e?��
�P�����
D�=�$̴߮}�kܑHG��*�����>��­�X:��鄏�׬�2�G�t�L�_B	� ���d�XO��n��5�f}��lK<�����#���nR?g��Φ���3m��N��1*?�n�eI�f�n���5KSp(Nx���o��}&�.��}�Ч��MG��̬+�~s� �� C�.�0�t�0�W����e��Nj��΍3�6;��ܟ���`�!UP-B���"�`NR����왏�n<�T'���sێ�&N��l ۣRķ��2\F/(�h|:�<����[�P�a��]|.D�-�o�H$%���JJo��2���4�r�>����z֦t������X��6�׉���H�d-ց�����@C�r�z�����^"nV��� ,	��y�ƎG�����r�G�`	,�F3�%�����]��h\��Bqڻ�7C>�