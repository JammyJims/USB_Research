XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G���>;��ֳx��j�i;�EXķ�B�(�{V�+�=jB���lt"�P������@�@�tq�����t"�^Ӗ�>� ֬�}��P�:Ri
4��e���2�N[%��(�E��OˎEK�R5l�✷R�yY�C'�
x�B�=Ń�T��8s�>>�ޟ��H�����C�H���`��<�o2i�+$ţ����*�z�މ���V`��v$��1�����hĄ{<�`�[o��86�W��W@ d�­��������	
X'�_����?��q��G� �6�6���tu�?�uےt�̽��m����c~��0K�W����I$�ޖ�u�Fuu�'�5��sY�=U�E���p�*��k�ln�bp}��6�5U�)��[�����KP0����"��������wrYPs�ڞ�l�'��|f��|�R�{��.I��k��r�*y�b�rQٶ��k�`Qre�+�L�7l,��$����g,����S.�:��:��bg����t8�O�=2;�5ذx��X�=A�4�p^Q���{�~?�pH�Ϡ�q�xC�� �����յWҺ�-	�!.g��N��b<�4�kQ� � �7K�[塱�k���e
 ��Z�)�y�Xp������
�\���n�y�Q��(^H\fS��Q����]=�#�_��+�se�מBW�y�b^7f>z�h��Z��T4�/>�S���P���7��j�B�%�I�v���@9�c���]��|3��r��*G�FXlxVHYEB    13ec     7a0���!ʽ��Kt��P��`��y5�,�S��d��������t�C/�q[��/vSWR�����NL�qI*nr݁70�+"����~[�[��׶޶�_/Sز)6
�<u���^��f/�?.�P��Q9�����X�7��J?����xHUF��6Y�|��F�3�,�]��SNS��B,mŇk��$���A��A��Ҏr�;�#h�Z�潃��~�x�'���zХC����;���4|�_�[{@���"E���|k��L������GW�YDx��J)-/S������$��� ��-��;��y6�������3�@�\��ՖAy����t|�I�	!��p���
V����%q�
��������ϨC�~��ץM��ZLȽW�܇(�!��6�ejKm�y�s���v��fB~C
$��&�ȝ4�_�u��X�}��4s=��D+������SϹ� �	{��(U�Ł�5Oc����q
IPj����1#J�@%���斞X΁�lZ~�?ߡ�S~�X��Q�5kn������O�mb+�*F��®���*������~ӻM�X�?�ɴ�$h�7��*��9L�d0�+� ��y�0�͟2�	�
��ʊ@ɇ�a�~v�(	ɡ��i��Иz��!}��
笣�v�MLH�����Ӱ�������V+s�h�k�_R��j�P36U�t�fF�O����aͺǃ܇�ۍ���Wg�i��޼9�	�v>�c(��A&4Q���ZƔ�6�ܠ+����zd�Hg�\���q�q��{۷��bj�`-x���x=�4��O�.�4�n�P�/ew�)�v�T&��`+��޳�TEԴ�pw�S,Ы���Bw��3�.L!U��j��q��(��Wס�#;xrT���Sc;�^D�!wR�(�*S)
�+DKր�Q��-��"��>+�<�&5�U<��K��'[��BA,qXR9��R[@m�g�}�Ḱ��mo�ɢY���+�_����d׻�q������E>�|7�I��a�+��0������p�OK��>}�C8�(v1����z��
�S+�eđ*�5_"�ٸ���ш���s�~�!q{m��1j1��\ }k�d�⭾��N���:���,��z�jP�,%�dցU�EX�#OR�}�k�5x�InM��th�To�+�3�]�`�����W˸"�YD"kQ
1�YG*����C�H�����S� Բ/V���\[��W�2�1hU�	hv���Ujo��]�}d%aF���#�@WՇ����EUdXz	ZC�����Xފ�����:s �����</kV��?���g*��	30��۞N~4K�5?ǿ�+|̃�R�-z�)�wG��8�^@
Lz�#)U���F��z
���b�GNf]�Ci}Ҧ$;�*k�&�K���w�i}�ݸф5MjÔxI�����RVC��rl~���83��>���/<�j����L-���j��_��̕���Ȯ��y��O6��k���<�f�w�veY�W�4�V�v���g��=/I��� Mz:����ؠx��~_!���2�η7�Ly�F\l��`3�cb��j����K��K,Im�!lG@,
G;�0�:�~hO�;�����W+�G�ݲ���7U�\,��ɪ}/�eC_�-�j8Xzd��Zo$�Lh��B��с.�9NU��X��x�J�#"c��_)���t� �e���F��a2B�o鳍0W�55����j�Bo9u�N�	(�R'�oaTڸ�-�8;v,�2�qԼпX6�9�����cy��w���[���.@�{�XAmY�`;��@�]EȨV����=*w��ek�&~`K�Z�F�}H�Ek�����h
b�{��L(E�ζV��ݖ��@3���O�DЩoqq�x��/�