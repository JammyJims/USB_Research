XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����dy A(7�i�5|èO#1L�K���Oj�ouz�)�t/eF���I4��Og�������a*b_?pm�o)j;G*Ʊ��i�<{�J{kZ%�ɫK�1B���cEl�WX���XI�\����KY�,f�Ǜ�1��4��Y�g�g���j�0�bQ+�2S:.�*틑?��ך
m�r�I�3X7a�Q��>@4�b[�����Ӵ_	���K�g�Cs�ө�\��P���3��q�_�瞕�L��S3���O�a�i"�ͭ"}Eײ��$�	��l�Lf���r�UkDTnI5��Q�wo�M(�[�n���f;��o\�9e�s���f݇  �S�ο݅y���v�����`����a���8�I`]���\�W��T�ג]����7gM�[����r�$����YX����)��k*��g��TQV88}��� (a�0@��q*���*�܆O|��*�X}4�\f�+��F��H����l�(�vsc����k�5��n�FUTYTwg��yv�RY��)���!8����o�v��2,O7�vK7]��Q��ER����u�I�����@�~�M��B�A�1�����I��v�Z]��K�/8e�xS�T���ʀ�(� -	PO@�T�k�`c4��{b��/?���JO�}�8��m����_�"�83��&���ʟMyk����E{���X�YuHꤙ��Yƚpfi*c*�dO�@�D�A!b=.i*�7\���6�Ʉw��i�|XlxVHYEB    2962     bf0�!z}�,V7dq�-9�6l�c�����o���My���(���ߩ�ZK�?:� D�	���F��� wR�*��%�@��İė�
��	��nf�e�, 1��T��x�_�i�8-�&�C= L�I=�k�z�w�ق��7@C&�R[�
�ƌi��<,�tj��Q��]���a��]�TI�U�����If��t;�Ӿ�跍���p�NM�,EMqq��<.-���'�ߊA8. ?'�����=�hFQ�q����߱�����Q�H�g��0�yI�5x��nK���]{W�]&M����/	T(�E4�'�^�%�x��ň4R-�)�ȴ�f%ԈV�*@jtZ�'�	9
���Zۇd#I]��c���0��[�O��ti
���ৱu�k�|.;�%!&��Ύ�P��hc��"f)�����T�B�c窌�V�:q
�#��M.���JҎu?��Y�P!�^��U9ď�"�� ?��ܷɔ*�iU���#
�u�׻Nӛ����09v ���/��L��})n^�Fݭ-e������Ut�MB=�01\�L�f�ꆸ[$w��ӵ=�8 zO��C�>�e�qA�ks���ܷ�Չ5�R�Q��wf�R�+ .����Y�Ѭ$�������ց/{a�>8�p.U7�m�� ^�DZ�UruZ��LM� �쫯.�k�{��; O#���sr�8Y�P���(F��Y����

��]���T�d��u{��ʜ�#qa ����`Y�E�RO��G�vD5�VQ�+Z:��b)*&�����/�+2��n�3��Fm�v\�"_0J���M��`x2oX�f�N��4� \�q�����z,�.�$�`��Wֿ�·u�.�}�[Y-H�� sv��� �m�Z/�=��_ ϯ��*�i�O�a�u1쏓Ǵ���^+��-�.U9�"�4�!~��:�
y	'֮��3B�⌭� ;{W�hܘ�cݸ*s���J����7���5��'�H엪��1!E� �8/}��Y��$ʡ��D@�Q��v��Zfz�F�D��n ���kT}*���PTm�,3��1���q��J�.6Z������~���E>=7f[���� ���>��������.�lZa[1�(�l�J:M��r��g�f��Zru�u����?oʪ�ϤK�-,Nl0X<��s�H���aN`"G��]�����j�N:�E'*�6�V+��
Zs��UּՆ!���8��m�K
s��S���lz����	���״SƉV�r״ݏ_7�	���,�)�W�^������ ��"�h��َ[-�B]D�Q�Q����0�KP�%�#�ն��+�*�=�T��r�zM!)H��L�����j}?H��ݪ�Y��[�����t8�)oB�0v�7������oz s�f����@,_Ǌ�;����i˪.�`є�j�52$�Zy,�q1���C��Y���V�t��ר���KLy�oӜ���#��[�����x�m��F["� z&$!m�]���b��W��%�,K��n�I�ߏ���!���!ݰ7�8��N�>���#k�ғ��p�P�O��G�>���� @.���+��ݕ�m:.K:{5��Jo3�R$��nɈh�z{ݒ�*��&�x��G�!�	���?�e��&���� F�S-(���u{ԎL�"���1GO[�[r�M
�-%^�[
��}FA+�č:��o�%�%Do��<|�{3+]l��g��fJ�����XZ~�5"�9�-iȢʩ,�d�'�*V,'���Q����6�U&��7>��x9m����1�1�L�[~�I�S�}���ys$ś]��S\,y&m�X`2.�Ԝ~v=9R�΂�w����tՑ
��Z-li���dԁz�aF��,�7����~�<�d���Ԑ_��W���a�u�\U�O��~:w�N�����[#��]�(�-s����D����V�1�����O��|v&;���~(���$��(��6�_j�o��e�!��@T6�1_Qd��g��Q{�%~�4d�l��R!i�T���h��A�*M�$��w��z/���{��w.A���%䀆b�X��oH���0`b6�{��\(�tjnX��0&���ZԜ�y�\�7"[�3{EuV1�9~�r�Me	�ˍ��Bkcz�|йI�ړ4�șj���sWI6��RBOkv��04��9Rܴԟ��T��z#x�%i|[��q�0�tRX��0��2���б��}�A�i�/�Oke(W�?���Pm���u�ʧN��G��n_���W���0�4�U��0Ê]*cϯ����mtl:@��'b�s��P�VH4�4�Epɺ�Yd���5�ς���a�C�ݢ	�X��ێ8!춑��Oٿ�U糁��tj��)��<���[xfр�H ���أ���w�WS� y՝h ��_�g��2&��K�8�H��a#b�5N-�mJa�@� ��w+�pNS!��ʘg̪hύ���;�����f�m:���?M����GR["b.@�*��j�b����f��������J?�鐱�c���{��#�b5��5�|T�'���$�S��������꧴uB�����tW�yQ�w	�2��h���K\c`<3@X.��j��c��SΩDx�*+<P���D--����ˤ�ZjV~�uK|�c�.\.�2�ɹ��7������J��sOm"\:�W����+�����G:�~M6��԰���Cl/��(�����_�3�"�cGw	�5�Y�Z���U���t�bdG̿�~�9i�2w������C^j8��J#��#h�6���J��ʂqh�����O�1J3'���i*���cB�K�ʚ�
�]Ue<3:�Ǫ��P8��;ގ��f/�{��@�A�0F��t���I��;���� �֧����[��+�@� l��8=�>��S�>�* f��_��2������ТG�=4ʀ�/I �N2�ķ�>�|�K��