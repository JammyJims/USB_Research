XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P9ѹ\�r�A���n�ܣ�!V�����@kd�>��7�f)Jw��ąwM�s��q��'	a�U��IB�/D�'n��%�p,0<섯,S�ꘂjC�?7S)�,�:��A7'T�$�������7,���T<}����S�l�L�,N,��1�K�ܯ�m�lE��}`u�֕��Q��]�-/��s��9%:c�"z�����R�U�a�h�5f�˸XVn_�[�2�]/�߁�;LW�D��1k��E�䧵mS�쿷��U��x�wVI�W�9�zЫNK��!�ma�R�{`r�s)�th������R���c���mŕvȞ!���|�=[�����f����V�_8�	$0�28�4�H�yg~��� Y���^�8Ѽ�ƞ3��oh�<4u��JaB��L�v�ݯ�ꊮzݬ@Z+��/��O��e+ii�z[�Vr4y�G�qeШ��и��
��r���}c�y��p��Ԁ��	����7�H*��G�>%Vk�h�'$�������W�{��;� (�t���\Mׯzv�X����hѭ$9;���2A�g�v��0ҭ�{.]<|)*�cA�	'EW��&�vT���[��K��ny�)Eh5���x��Ҩ��H������6��Cu_!��o?�/뤪���@�9s�Re��U$
N��@N�,غ�Rұ�o�W؁oL�\NSU�2L�H�� {��H�=kC~#���=�/StN����00�w/�ͅv����a��랺���	;)%�Ztec��XlxVHYEB    fa00    32403@ǧ��پ�>�����䃪�H�����a9hiL�#'��~���gS=�ǚ�2����B����\��~�ʹ񥽍
ވ�w������V��eU�m��!������I���\Q�}aj>G��hV����w�V|�бGc˞�%�-V�	͌Vk���[�{0$���V'?�"���`eR�ԹSw
8��N�u�a�5�}%��`�Z��������/��!r�m��c��uG�!������%d���?�6���h��¶J�������W0U��U���-݈?�݄��&�t�/t-��~���l7@1]C���a��,�U��5��wDR.7"A�M�y��F���g���-<����L�Og�#.�3�?j��u��~��2�L@.��5��*�#��Xs��0�l� OˆH�|>�ޓ(��y檠 �n=�i`��+rź�=�|��2P�'0���o꧵�l	�Aޗ��(����׍�W_�)m�� ����2ԙ�R�[��/7��=�V,���El�#;Ɠ�o�?
3��Տ^���<Q�K���};�g���} t��2)f�l�Q5$�}0ӈz���ۊAϯ~R3�Mg�[3�O��i#9�����O%�I���]c|e�f�E��D:�Ty�GI��n��8�X��Q��qH�#O�����=J��-E&욈��8lˣ��|~��O�}��ڽ���u�n`������v=�)W?����D0,`��	7�;LO���BE�����9�`u�Ţq%����>G�	�޻hҍ��6���5V6�srJ&�e���b�g$[;'zG�"��� � g�� X�ɻJR�E�BwD�f{��+�d��of�_&$��y~<�0�y���s3�kv�O�w�%!���V�`���� ����)({ȫgu_�*��B�0����8�Gqj�Y� p�m���kq�ܢ(�_Y*�v�|l��b�X�h��G	_��A���od�lZF�%�s����]^�h[���Ҷ��/\ w]�`^{yn�QK���T�L�k�T������﮷���We�y����"c#��\�(�M>��5}��Ї�M̈́�B�'*Ū GV�>BS{���ɏVk8���gwO�S^�ϸX�zHv�t���=}�Z 4�R���DBYs;�.���(���E.����ZUNj��4+����d%Ⲃ���^�(~������3M�����(��P��.B-\R�!Y����n�3^�u����`גH}A9��7��U�Hl�q��'+��S0�&��|a�c��Vk|�{��p,��Q�5t[�
��ի �쨣��׳�1�"�J��lp��
H�������J���Ȁs�UKr��%2���U��>}Ѷ�郟sVP�Ŗj�<��r��-��IJ�l�Ys.4d�A�T�HY�j�f%�{/:9c�v#{:�v��lYr�z� �A�ÛTo�R�$`B":ڎ�mv׸ �1�wg��԰���Z�a�" ����Gܻ�Hq)���"Zd�fln���'O���{&���A��z�By��Ѳ��y9b�ȹ{CdY��Է%�]o��*n���:��LO��Z�ZU;�*|"'󡬂KtA�ƴx��4�;̃�dgK��%Z�&S �+�Rj���oP�j}�ubS���:yDwC+֋���t��O;W&�y��x9���ׁ�\g���7)�}��JP��gג̵��5�Pb��_��Oj�O��n#�ؾ�����cc+̐��pӘ�R�/=ϔ�M�tY��ޅ�A��K������&��+�X�P\�5��`t��C�=\�[JHX� Ru1Q(�ڗ�Z�Wb�$f�"Uy>�)}p'���38,��OAX�G�em��|.;������A����Pt��Ֆ�f��q�P,��t�
�.���J�9�7=�+�C$ote����*y��6u.���;�AM`#�z;Ĉ2~�3E��w���K��4D�<��2Ϻ����3��z�"�i5�1�v�>*�O$e�ň;��dK���m-��V�j5���#�	E�ǩsL�"�+'	2v��$1��f{���dS��**���I�-�|��K�f����e���JL���0gu�z��[N����U��DX�'�¹��"	���w���g�_�ް/���R{����E:����)q�^���g,�Ŗ���=���	�jf	E�"���Z���.��Η���Ht�%?�V���[���iU9#ʈ��<�����i����h����]wq���ݽx�|r�i�������h�y��\m챇�O}����#`bG!h�?��Z�Db��4�w���-�C��m�i�b� yB�d>/�N���6+eh�7��"cOj�p�ck팛����ea�`)u=�w9@��T� ~�"�.v&2Q���~q{���n�p(���r~�>!o��|�4PnE_e��2��9�/�����f�2x����y�@(qu�FnG�tV��x�H2��)��h�A��o���N���Cj�.L0������k��E�pG4_��m:���ˢZ O��h��A+#�8�C3B,���z���g-��"��*oDV��R}3�����Ae�o�*�L�#����!`���3�aU'��j;>"�����YM�x�^
���c���A\��nL���H�<�>�L%8hnz��;X�l���CO�! ��2����H�6�b^bRq���[��"v�3Yw���!=�m�Ɂ�=��*���9�L��X�6 �c���b��R�gG~�4�qu��#��(j��N�,�!�&$K�����$��U�2'�h�u��	�[����m�j�)�Ѓ���D*���(�-]��Y΋{���y����9t��]�9�|���׆�W�0c���~Ɛ���.��Kq�10]M��y��l�z��L�-(������H�YT��c���e����]S-�a���	�6��
	�b�ܹl�����5���ڒ��n}�7��3/i�X!���?Ml_Ek}6�@C�)9�V�؂�>d��Ui�mj��6��[H��#��lT$zY���JHÀ�j^���(5�5T�s��%o��p�d;�����}�8;�����BG,��S�w�+smP�%<�ni�3Fjxg�lƞ�
���^tuH������Qf���C�:��3���{,4�'����[�!�lO���gx�q�����T~3B���ȼ��W=8������w�k<*���$1]I������Wo }^h��6��t��Ҟ���Rd��ȴ���j[7I��Ic�{����vQ���� AKI���ˣQp0���+^.�L�>���3�A��忶����"IzF���.`�s}��ﶣMWUM�k��"\�1I�E��3Aҽ�i��1 $��E~��$�����::�w�>?�0q�♅-_)ӎ�p0����#��x�F�L�	���0�c�geo��!�\�ӑ	�P��#n��!�Q�e�8U�i"��Ý,f-�I۵��{�J�O�喁�����2!S��fj��0����y���%�v��1��K��YI���'���({��������)��]�����1D�sm�q]����W�v�̽y}�B�T�vB��_G
�y�F�?�J�ic�cD&(�4,�n&W��؇�5r۱Hi���w4�ҟ�r�3�T�_3'��!�]l���f[ j��\A���|_9���d"��PJY�Dl��2�E��j�;*��ӌw<�В	� �y.��Q�LP�	8G����rk�� .�m�NCB��%�|<I�)��@}��i%Ӝ_��c�6ǀ$���S+b�`�#�2E�BsZ��]�(>MCB�`g�ǧ'��9ͫn*o�9G�}�Zq�R���d�_W[�@@%�)�d��/�V��X��VK7|�7a�$r{W*�ͅE4ߋh�Βç�]@ܙ�"Mgz�����Хa�Mv�0���k������1�.u(�2�����'���xN�d �F�:`crD������Hŀ�t�	 �2�"���A�))ޛ���v������G)@W����^�ʀ��xY���aQG@���k�� �o�,�|E$��T{ 4XV�F�dz��@����i����%�.�t��䚰�\�אB�!�e���x����_��e$ۜ^������&5���|�$�0y��<��Od�M�@z�������X�14CI3�a9��&;�M��-�
9N�G� �|.��6���:T�������l��^Ǻ9/ϑ�3�K��+0t%Ms���!34'�����,���*��A7�&OH*<�BTz��}�O���8��G��­�t�d}���;H�{BS�1� ,�W��s*ZZ�M�Cǂ6�&,�P�}͏{���"m��żt�_.(��f���nMJBփw��<��Aܥ�	X�!ۀ�u�/�9y���r
���
NcM5�l*�S�z���ҟj0����|�c[Y��-�f.p�]��i��v��:�)�D���i5m�)��w�8�A�E�'�d H.k�0iW�c}�bn�����¨�2#&.�g�Eǚ����Y���d����%�� �f�c8�٨N��O�I�	�x�㰝�:W{y��]�~�v&�;��r����68M䀫��8$O�q&��B>�l��͍��̊재 �t�8,�ݥN����d�L͆�l�Z1�LsA?�,�Ɉ�Ë�j�O��d�t&�;�n�C��W�]���xn?��}U��/q��jn���㐤�>���P��6��� ��\�[Pj6�Ef��p�TV��ۑR����D1#Eֆ���Ғ���Ec�	�hh:!�ڎ/�04�+�ES��-[�E����+��D�� û�􀜅��
d��D���@ux*�~��L�\�{�d��j4�#�'#�*�5�LSeЦē�s���8b0�*g��J��B�6S��_CJ�ly�x�{�B�`��g��xOU�h��D������$|����v�啟ms-��6��	f�מ��7�M�O@S؅8P����ٕ���7�0�s�N;�����O�='K��rXV�7t�������nՑ�D4�����)��,�.š���聢䉟�<N�〤L(:v���������)<�Ԧ�P�%������?<�QY.�Dﺚ��	���k��?F�n���J�B7��j�ٱ+l�x(�ݲ�Z��n�)[|��i2m�sA^rd;��5σ7qq�x�R�m����34��2U���7��<)h,�s�6d?�����C��P�$��rs�j���c�`�ha$u�~�1�hے��;��~���)��G]I��v��N���NL���P�a�}�x��4�Yw��M9{@#�T��c�IΩ�@��z�8�>2,V��K'N�����(��7�b���f$Mt�O����'��
�d Z ��l�7�y�4�~���gĿa�Uu 8yV.�lQD}s��4����dFC
t�r�P���3�T�ù0�6����J1z��<���>6��2�H��p�t�? ��5���-=d�2��Z���"TXz����A?��-�H]�R�4:�s�9�}��B�B�gx�]�X�J>4IԌR��@���� ҋ]�RdY� 
�Dfr6MZK��֍�m����2~p����d9~����tn�Kt7!�S:];�ߡ6^�
6n\ر��N쌞���bf�w p봇����x���o��-��nL��2�����O�:$��T�G@��:{�0mѲ,��>)�FaΧ��i��=��F�i���Xt2�Ĺ�b��h\蛻�U��y�!�4��.���dG��޽l���G1(�8����'8o�zB	�dN�VF�-� �Ԧ����Xy���&Vr7j7���w�{g]a��v�`ݑ�h��8 ���(�����+h�O�璲N*|���Q4���ݑU ���s�2�ѷf��2]^�Ó�C��{�G���=��*Y�^�A�������?_K�5�B�A݀��F!��� ��#GҾ���m���rW8�^͘�)�'-�N9�f/�6&C*��aɓ=_`y9i[#+�Ö� ZIt�A���K�}�.7)*�6�iy��b��P9/@��<�l�B��e�P3;�\��.|
<�q[�3�W�sv�:����#�]S��_�ڡO��~usS��'�k�%IX(�賩�/S�'�����q�z5�ۍj�Lg�Ss�c���~�@��c�w3Z���ՂLn��U��3�m
���O�����������k�a�M�^���P���eW3���$�2��[@_�?P�>�E9�hx��O�}9�+-8��0CE�U��Ɍ�1ގno�&&�X'I�DJ�*@]mT��'��J4%��a.����ǔ.6����C��軷�,���_ 錛i��R�6c�/�o~��԰-�'zO�d.�.�k�{נ��_ W�ևyW�u�B�@c"��q坼�	^J�W�!Y�� ��,.&��~�<,��~Γ�=��"�=.��x>��@�YH2��'����V\�u ���ƶr~�c*0׉%*R*xN1f��JE[�g�p�:��wF�f�ʭ:��MK��ٱsZߐ2ƻU�w8Z��oDs]��`[ŗ*�󐨭�p{L?y�U����,={�$��bL�w�pL6��"�.�R�>c�G�|0�؟�.HK'S�"�o���[f-�5
�C��?���S��2����7�Ğ�Dŀ��g�VM!�n|@B��Si$X��}U;��zˆ2�@���BPM�}P�hX�d�^�ا.aE�M��EAٓ�S���d�+��z�W#*:�Pͭ> J.�gE���f#̦6�L[�?�	ι9: rS����^���L�I}X^��ķ�++������}M�K��9L�g��1C=�ʅ �s�K��?5�?ߛ������oѨ�&�M�1�v_i�%�r,7�Ph���J�½�N5����Tz)�Ԩ���|��~���2.`n���7����sI4q���*���P�ǲ��3r�G�k�tX�h?����T�]�|)����Д���"S���pq�@ېeG�2������%	v:~� D	>���-Z�m�jB.�r�u�՝��ͅ#	i)7�f��\2�%D�֑���۟�a��
�@}Y�?��@�;.�B���J�X�M�No`L���x�ŀ/	͗׈���A�K�AhD�#첽R�T�|@�*�&4����D�ˆ����G�g�ƑM6i��]�����c1��;*�X�>;,+�dޤw/����|4G�1ь�v)����4G����*�Ͳ�7�B䶒G�O�:��ֵ��a�U��>��5��Z�Zc�6<�RX �����7��`q�ቬM�UV�K�w>����48c���U���! 8z�D&�?���Pob��б�P����^��e�k��~�Ϯ���Nߵ�ѓuz�q7,��|�3�!/GQ6W���\~<>N|�(�d�ީ,E��@N�󊍡>��.��"� �~�`���d�[�D�\TU�B�N�V� ���ρ#�H���faڰ�M��K� �����p���} �&��9H�W�9u $޻����Q�����nzhg��
���g:8
�Z�/�H�6���������KƝ-�S_��C��%8��<��:��i��z��y��hG����2���)���raJT�x��"z���+L`��y�]����ϊ5i��{p�l�2�����T���Fx��{��d��"�_Db�Ş9<�?6��e�g;^Uw����Z.l5h�{�,�X/��t��`+'����y����.��ݕ��$<�s�,g��,OsH�5��6o*�Wî�?1͢>�2Wh҇@H�����g��6(H&$#`�Љ�d�ue_D�%E�QA�Ù
7b�p�-�d����Qr�;<�����V�+��+���)!��Yz�뤯)�'��9۹
�ǣ�� �UЀLʎ;~�Ƌ4�{�*z��ZC�>�/�<�/�~��h�ɐ,6�փp�����OL����)@&�me����%�	�b8`�f���	�o#i|ze֎�g�J��L�z$
TRT��>�:����#Mqj����� J�+׷��~{��P �`>c`*����#������q,5E=�����Eq'���b����Qq~ڸ!#CT̐�����ܝ�����ʽ�c�b�,�fT�H�#B޶8z�lk��N&V�L��,�z��DGyL��9gC�z�Y�l�f���,f�����Dr�_��?�j�+9OP��rV�F��{�� �\��P�Z�F�r��c�oфq���iJ��v�R��ʙ����?��T�ŎP��Q�n���8�@�� ���հ�m���k�V2KX��9=��"h��Y�ﲾ<u��\-�KL�H`;;�hl(��̶К�՜t��!�{�x�Z�G-A�kJ�Io(���h}�1��G�K�S��@y�ś<�[���U]�6�~@�u�]�#C�mm��e���f�Qm;w�x���� ���R�8pӂ_����>(��������l;oaT��u<Y��Y]�+�){�17`#k!��̛n�W���������B�#��\��kvX�-^��-^��+ h�+^$�F�+~4��{����
Z����F �<�o�Ѩ�=e�W�M�i���<�$q$y�U3�-H��H�q�?��/o��H2!ܳ���$�t="���7�d����`
郷��ۿ�g�5�S�~��~�4%k��1d�-�A%*8U�L�i,$]0�
"�����Y���#�AU��=�T��?o�rQJKxj8!� �p�_� �)R?T3��K�����a,��ǜ"W���,��lk��pt%uYJ���Y}��p
��$+Ő7�WI�@�+�ay��Y�����5���ɭ��jSK}˹�_�rZW���Z�N�!~���d�s^mxXw�������ji��y��(W�ӄ�~�	�,�]&�t����B��
���g�x$�g4�+M�{�ҋ�ɝ����VC�]� ��c�<��T�Њ�d�ѵ�ʻ��� �r+F�=7�Qf6B)��)�um<VF�����P�\���_~��0��I��j4��i�D6�y]�xnL����}+͆ûKc����щ]�#z}��qr�� ��a:�1DkȒ�mu<��qK���Q9��9��R��)�7�+�i����4��:UE5GjF���y��FB�7�7��YR�-.���ז��'�Aэ`�1�!�G���T�荜Ά��$42������)E���V�}�!���_�J�h,��O�R+*Q:0u���N��-��@/��I ��A���8�a��Of��0��`�(�N/Y=�w��J/�9�Z�e�����P�M&
�2�$��c���o��[���b $��՝v)��=�¾����p�F�̅�qm�t�/}D�)������s4K�{�͊��g�>K)��ѱ����%)�
�J��)��@�pnk_�hH>^�z0�-ۈ/�#�W��������I��ԭ_�W��^���;�8R��2E	���q�y��CJ�w��<����O$�z���*����I�Ր!�rVU��Y��9�$�-&s�v~+����Ҹ����J*0�g����A�w��G�Ǥ3�-��G�ʸj!�H�t�T���l� |����y�U�W)S���@v��N���&��*��t�,�X�� 1����#q�j��u�.�T�I(!f�~4Ũ�Ҷ9+<(c��o߄�x���p�-5�)\�<\�u��=ٴ��q�Oǌ�X5�7O�����@���X�_ÔJ��C\g�|����Bo��u,\Bn����ezZ$��$V���c�0�C������g���)���M���$���m�տ��m��Bͨ�!�ަG�� JW	��y����ԬP�����Ϗ_����4h:M{�9^�ղ�~��n����=�r���R���n�B�l�|���2on%-[����<Q^����3юe*��A�1J�ü�/�����}~��ɑ"��8����u���Q�������C��SP<2����7�����ѻ����j���u d8~�˲1�CJ�f���u���wX�o��mM�5�������[���U�6�:a9������ap	H_"�nGN���t�}{��_8.�7�b��s�o[Y��c�!�{8��ꠦ�F����)�
��m�K@n1p��d2�LM��!���%�怼���$�2kFi�e�G��Rq�M��Dՠ
�OP�b�\�I�p?	�Q �*;	ADw{�C�oB�����̛e%��E�I����"��B)�11;�+:.c��s`�H��d+%��GՀ=���1��!I�׌��V@���}������|PJy�m��[=�@Qt�E1��W�߁��gc�z�]-�_ģ�ʐ�&K[��,R�t�)�Zf��C�4��4�ӑ�$��3����^ڻ��S@�=��f�A�r+�#d4��UW5<��j�c
�7:�y~����1NN	�>�Il�a�E=��tԡrL�nS`��B}\�[�<����Ik�`[}U>��ȤM�2&��E�ۘ�����6�x��I�5W?X���"���>�����#��Zj�o���.��'��"_څ�F�@�K%@����'��/Z���sª+C0����Y����B~
jFP�%7�8e,�B� $^~^���<�惸�ђ�Ŏ�+�]}+�v��t�Z��_��c.u�x������k6Y���H�B�����Z�6VO��3��"����*Ø|?rx�T`�����"�'p�9����*�O]�ɖ��a���?d(����Nz� a����L���AN��
��T�pŶ����f�V#�'�d|�Kl�X�Vw��E��ί��И,�wq׈;)����mG�C�6lmj��Z�)�� ���tv�J��n_2єO�6�I�����Sp]+)%��
$ĢcT�J4tn��=��^Ċ��R���ֈp�����d~�ֳ9U���$���Q��I⒩GC�S;Y�@�V/�|ۂ�;!����^R&�bMX��f���7����7�)/�1Jd�#~��856[l�5�,����2��9���y�8�g�STwM.�Ϳ��RR?>����{Nh���f'��t��)"KL�|8���[�GQz��ad�t�ۦ�Ƙ���� &�pU�t�)��U"�0t���o̦� �d����ҁ@�n�<���qUXԈ�ǌ���ivШ!�x�J*�V�j��!,�4lg>�w���0��j"R��x:~�4��߲2 ތZf�U�>��I�����F��	Va��K�%�A�ht�w×&�y�G`ƈ'��'�(����7���cץ�E�jâ\1}�:��!> �U0Kk/(�۩r������#E�iڲ��'ҧ���W�
��7Y]!ᬢ�T��;�?Q���8�멡�
����'G���~7�*�ϫޖL��
#�	��Q�5���HK�~*�$��d5lJ�&�K�
�'����.1|O�Ĥ �M��x�e.���U:��A�Q�������:hހz�#��*��eym3���bC�*X
�[���-���K�ʠJ��O�Yt(�dx�T��*�Aů���Vpo�N���"����Ј=g�]�:}�F�
߉q��h�X��|>�lo��X�o	RT���5.T��6�����q{���1�p���t�?�]�gs#�Q�-��� 7Bɫ�x:5]r�A�&U�`��c�������&>�B��VoR(����&;���+�K^��0�b2� iC��n�E��;�}�y�R��ZeiL��,_*�I�	[�E��	�렽�|�ۓ��Q]����J�]�?�[�P̙≪��}�-�sj��"�mU�C���h���8 �w���Зv��sR�3f���𜯂^tc;y���$� ��Zԫ�ppO��lSQ�ִ�@�2V�N�t b-8bLNՎ�����wG��4�̱�F�& �ASK�I!��]9l�)ٽ��P.�>�,5�Lk��s����=��n\;����pڒm.-G��)�j��[H�	�h��E�!�Z�=�v�\}�a3�U��� ��=^��ΖT�ͧ��f�H��^%�o\��{�ܐ�R���� ����u#��i�$�Z�Ո�,E	�\�%��5�^��罍S۵�t_B�C���'F������=i��1�Zg) 2��Q��	�)vs�B Z��xg;����$�n\��:���K��q� �!di���v=�?��8L;��΄ol=:"52�`�n�X� ��>I�d��K¾�'�!qL �5�z1�[B�,E���%��'��\(~G���m�u�M��[&��mH�	��:A2G�)���Ԃ��t�]�^@��(H�����ݐ3N	&?�����8��3I� L��@���b�7Y{�j��!��4�"������/��CG�h	�"�hc͘sx��4�1=#�hvS��.��!#A-��"�x�@Y�u��j3�6 f�?��_��"^{̑��WS�������L�WN����{�(5�Y�J�v��$���\m�����h�A��ӻ����[�I��r�a;ՄU�_{���\'�0�ѝ���"���n��v-m�1(뒘�XlxVHYEB    b2c8    1cc0^�yj��H��T�F�?e��rD��ƀ<;�d'�±���ɵ�Yдγ����H�R��$��3�E�<���Dj��=��<�קӧ��Ę�_�]>��/����j�0TRU;·o: W�����bm2�RoG�i���W�Jq�������u*8[I�'p�%Iv'c���EkP#���Ę|9���;���E�(�!b6�r�^"%�
:��<�B����N	���k���
#��[:���MV:/f�'meY�q�V�Go��{gF�h�z��$!i�=�"&�h4�g���&55v/ưu!�V���f$�J�N*~u��!RS��a:��p�Ӥ���rO;���g�Ä�ϑ��6��ƪ"ԇ]��Q��($e���O�Yu@4J&ǛԒy&�_03sD�=�O�h��t���ح>��!�&B���I�n��{4^���Ƈ��*'�Ü��!�=pJ���ar+���
v���{m�c�,����g2��;i/���:��Wݧ���;A��_�h~k�?]�;����y�+��0~�� z2ec{8@�ΰu���@��G��WmD��4��ҭ֫x!�-������1ԨB�*�@����XDz��&@��j]8��S�gX���
���k�ē��ωW���^�S�Q�	n�߂4�K�PG�v����3�����̧�>p�����$0Ը�P>B�����cw�l'�eqϢ��D-��{[��������o�{�顎���R9p�)�rO��ύ�.�d��HeD���C�r7�eu.�Fr޶�裖�={`����p��Z�v;Ƶ��䜬��Л�d�-]���vh�N8{�A�̢l�}R�-�U��,��N�axV�=���)k��1���������ɱ���g *زE�<\2��!Jxs6^U|����م�&�ҬI}dw�	��;g���P���и�ҡ+��q9,�|��M�}B��&�A�'��2�.1v3�]W�9r��f�+�RS%2i�/�
�Z��_gp��������5�� l��Z��B��'�nF���JCC�?+�1�m�����J)�-N[�6Ol`�3ǵ�s��)	�v�oP���Fg.ͮ 0�G_Qg�Чv.r��]4	^��+0���21ØC䫤sk+T�9��ϲm/����]��D�Ȑ/����a��H�i�ʘ�,�7ỵ]�\��XT) ���v���AX�}ju������G%�Fk���1G�����GAE���sA���##OR�ҏ�(<P`���ln� ���v{)F!�^4��`EĽ@"��<��
h'ÒI]�=�X�s&�3 ��p�>���;���é=[��z��7�:d�FĨ��ik�d\���R�r�,�	O�r堡�`�=�'La>AvV04,<��˗a;�[<�W�t0NjM��"��p#���E�'�}�
�W�L��&!�t�I�>o�����J�A,�ҁ�µ��o�
�_���}���"�^Src��O-�������T����)���C�b����I��+ȡ�X'��d�K�����%�2�̓%�ey�#��վ���s'MJh���Z��"v�,���0|�a^?�:]�e[T��-h�"��&/f��a�F�����K��86�dǻt5^����'m�e!+Q�QR�S���w��VF�C�'I��n��+���z��H��	'֏\)A�����@سD4���R�%p^�_�&ʐX�e;�2l.��,٧��9�Va0�kЉ9�J�!�a�TJkeM�(�ߘ����l��s�x^��:� Y%M����J���5٣k���l~�m�j�[����z.�����(�KC��'��8劤�{�p�7�^�O>;�W=Y�r���C�{��M���X�k��j��'���`�����_2hǆ�v��+Q�H�42'u1�m��Ϳ^�v�4q,�SeI�y'|��)zsU��C\�W L��	&�;��t�mY�@�b�YJ�AEE�ׇ^�)�m��[�J}���^����kթA�z7���,N���L	�u�sg���V_�=��c=C(�'@���zva�x~��:�`G��l:�U����k1�|��;���n�w<�y�yOV�����a�|*�����������ac�"�Ш��!�C���ej��%1��V��gq+j��,����(��|h-��k���wDˤF/'����0�GB��C�-�L�JyL�#�I�*�4�E�J�/?09V���K�A����l�ma�EAU>y&���P ^�ښ�%���8��
y�Bà�53�P�o��}��|1G�� ���l,�����|����ѫ6w�{&����eozO��c.�N,�\0~U�S�$/&W�f����b��G��(�DXn��C��D9�Վ1q[C}��sO
�h��y�N ހ�d�d;&Ԏ��������J�0�F3�HȠd��������FS���9�i�8��{\�D����c��$}c�+�8fL�G[qʥ�x���x��m���Q[]թS��]�.���'s
�Gyd�<4�Uy�R4�3q�v� ��B|�*�L��H~
�:Z�o�=Pa�YH������L�	�,}*/EȩJ~��H�s~�Ahw�Z�~�HB�½�k�m��fm�ou�b�Q2J�k֒	%��j��ޏ'�J���h�2+�P �?�q�C2/U�����Q���I|�9?P
������V�ct^��J9��EnQ3����k�K�����g��"�y(2���?<{�yS�D�$k���]����)��/X?`�I3yz��]\����B�s�lek�q���5��e��s�n�F-��Y���Z��*�F���{��F#�
�E�z�QV*8�I2�[��\��'���`g�]a(:�Tw�;�Pu3qLh�IR?-�޷����do�!Q�j[�3��ý��e�2�%��Uu?(���7�>a;�� ���}i,EO��E&IR�d3}��Lq�%�\a�$��
�5iK�8��bl;��&��o{̲����;B��LK���r��Ed����210ݡ�����n��&:���;��u��!_�#8"�Cj8�(+�ߦ�5�oz{�L�c^�'~y܋W�oh�0�aU������cw-8¹t�qe�R-$_�N����[9��:��u�0�\ �t�6@sݒoXy�|���H6�2������5��0�4!~�w��[ѾT���w���S#�j�&��QOδ����dT�n�|Ls�={#Z�D���ۆ} l�_��,���-�d(��<�D"U�z��U���ԊW6�å�ȧ�3M~R<�E���/�My�,g��S�����<$ѽ�I�Q
FVCH5�+�#�]j����%uQ��$ӈ��>(����#c�XJ�(jR���E��5^U�$�����f*���������m������v�8�{�H&*�3���zT�
"��?�ƻK��<$�._�{�줨U٬tC�k!i����?�/9O�^�U�� i��Om�G���k����;'e�p(��Ƽ� X1gs�����!���k��fSpk�c��X�R?���E�%�:���lh��W����es��R�:�2�tK��O��(#��� MiSH���6��E��Kn�2��� �A��@L+�,RĨ�:��(����p,(m䗣H�Wtwn����˓$,1W67�@�p�[U�E��s�x�vi���!D��I栂���R��J�5r���u�+� 3�?������k��/6C(���_/KN����~,\N�)�%�R�*�R9��=��غ��|�;Q�K{%��dk����h��P�T\�D�S�z�����# H1��4�꾐Hp��v��1Y���d�g6���i�)�ȂP?�������ښ�U�.\�?�
�W���隷
0w�8L|,�s����Ɠ�"��?�+��p��{�A؛&�A���:<1�k��H#�� =���m#�����+d8�a�l�����v�\�e� =覘���sR�b�.c��J�t���;3�7��� ���F���v8jc���T� �3q�F��*������x�᪦���P���!��d�j�)�L�� ��L%�6�9v.��.�>��U]{�-g~��|)��������X78�yVg�"��Pl�$AF����IljG�p+����0�s�/Y�J��g�F��HK�t����@��{aC��.���E5m)v�FsrR���NHYM�ֆW�W�B�� 3ՐF��d���F�$6+�j�(��U��\1Q��:��M�O-�#���Yu��(6h�>%�Yi%Vs��$9�(80��_�Ѵ��Յ�o�D(�Y�wt�✺	w� 8�>}�ri>��c����}�8r�м���m?R")n+�2������w;��{����eg?�Jz��Qe������[�bCȫ���R=A��i��W�k2¡b!�s��w���_�>��z�e�k��n�������I�.��Չ�3�.�eP[��?>?~��n��@7J�ł�g�]E�"�3�{��`�p4,'v�mQ���%9����)b����[�,$���<����H����I��i�+��mW"�?!��}�~��.������EY:�~{Z�Eޟ��� �1:m�b�t��o����Yqп3V��p)���$��w2����(o�%�D�����a����M��*�X ��35g��IҨ9�ͣ�AIZ:�.00�E�;/a�/�nMs�;ި&��؍=�#��Q��_"|W�/�p��F�`�:�5�Uo�K�i�ղ���j�b?�尛:�*��i+ٜ�;WTH�9�c~r��C�$BG��'��d�r7��>�l��=f�8wԄ�1H����z�i��8ЕE��lE��NJ��/����K�o�e���x1��o_���&૤,��b0.���h���.�u��l+/ou�tJ?M��@c[U���_ՠ��ڥãH��m��_�Վ6�ӝi��dο�mw�#	��J��8���"uE9t�NYJ~����U��a �0B.�E����y�G8p���/��S�f�%���s^m!��*��,)�}p��傪��%�_fǕ~j����ൃzg'��:�T_�0��
VY�d����7�Dn��Q���0���ڭ�t�*e�?m�ݪ�a�{�H
L�����r���0��&Y ���"A���?8�^�>/E�;��7!Z��h�k���q�j]z���2��X���茜��`�������7#���;��rYk� ��IX������>O.z�JunӑŘ	�����3�ڦ��M�ľ���\k�����`�Œ{HM�ʗ���TT�ٖ�$��)���I"?r�G���_ʢ�����3�		��g��֙������l�ˌB{>U�� ,�4v��O��P�-W0�H�'�-ǌΠY�$��t�l�.%{/'�����(F���ve>@��n`� ��{��׈A��:�Q�L���y����\w����� 9C��N��2����dq2���`���s���_dG��;��Q��<��>D���u�L|�~�.nG��&�f
	��e�Oئ[ҏ-�HKr0�
>��,���ғ��[4n�Y�5�9!$?��ڮ���g�eA޾2�t�ŝ�J݆������/�\�uE�R=�/�c?�g��5�Sr�H�mS����]yb&)�e�EYf�)K|
�੯�gy�{�;�CsVԱ����	C�/�q�C+�?�Fe��]�T���	��պFzZ��1@ӕ��W�b��TɎ�>ea�����E�4�1g���T�(��.������ تp "\;;{f�b����x�NYm�Ћ�����T5�ʊnFj���9l=fp��>�3ӌ���� ���X�Qz�s��.�{c������B/�e���V��i! z��1}�DT�KI'uL|[�XG'�w~2;���Q��ϱ��Z��it=bz�.j�~�ۄ˟�l&����í��@��hF�s��~DU�1�t�I�Wg�ʉ��<u��q٣ɇ���k�哊k�Y��{z x�9�����t%Z#����׭V�#��_�*�c� D)V�R�=����'07w��y�U�(A�Q�6�ׂG۷�1�H�y.�o���J65V!t�*^��T,\��>0:�_!��,a�$�s�T��~7�|���5���ZMx�;���1h˨��Yh����hB1��tQ�%��G"�.�Zf:��RV�=�
So�����qR� �_����h&^f��P�0E���Ϻ�T����2�tvZlf�6J�0��(&v�=�;�gnFh�Ef=��ʲ%��9�u�����y�aD:��C�6�	|�ʟiX7��cV
KA�?+�˂��e�M���U+{�{ lx �����bl��b���,�'d��!"5��V�G�Yi�/�_�O���T�Q�|��,�~�3�Hst�?��a��-y/ۂ�}H���G�"kT�f.�/z)�w�c�c�.bc��d}�^c�9
��U�I�T��a�Ԣ=5�5Bd�m�j�~E�Rm�&���~hx������SY�V�h�r��?�73�������cy8ĉ�?����K�ԫ��ܚB�"J����נ�vy�R��|gy���Z�M�~�qW\��C��������]�=w�}Y'�� ��$���iy4�����1�<W�U���T:�W�h���C�Ҩ�-�cUk!�qGݮ�ñ6�WH��S�
�RpB����iH���&�@�;��S�����)��u_=5�-<~�t\�n\�)�;M�������F���%�J�M/�7�*��+'Q�8s�Ya �{�J�C����W�����"�L�M��b�!ecJ���||��>�����3'j�>��)�fwI�k���Sb�)K��8b�$6�n���!`�Zs��穻��2�3\��5�r�x�~>T�zf��$��	+�&v��j�5��+�3���!�kC
W�X}�E���*�|KXezFiT�r{9�Q����y�ȥ��f��t�E�Q��:�W��Q�:d����t^+o4���?hy�u��𡶮�T� iY�^H#����\���������V���H��>h���'m���q��ߢΥ�&�a���q3�ч��LY�W�c�@l~�w����RDS�<�t�r���X"ֈB,������xvt!H*�`ؘzI*q���<kHk�m#���qh