XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u��ر�ty�1�˘��=�4��W��j��z�(.�Xo�W$��y��ǡ6��z�nl��}M��O�b�����A�N��P��[��1Q���Ύ�.�w��vu�,�e�-��4���V�Y��H�����#�"�&��� X��#D�BdN�B�ɭ
�%_��陵�<#���m�y�9�־y��#R�B��o2����L�Ǖ��$�-�}'�v�+U�*���C�Rh��9�N��^�����!w�����2y�P�����.�L��v[��|�c���qM�C{�\o.<��n���Eܨ����X(�Q�B�Y>��R{o:Ekdty]WN�B#���YhG�0B�=�P�ߌ�$���m=�VE���M�ٖi��b5㕎��� ,V8Ȩ����A�T'X&��)��ﶣ������)񉂀Q��*I�҇>Q]J$ �����N��F���S��p�ƞ(���l���y������,g����I9`�/�0�<�����'�4�.�V��:��b��n�e8�fαl*p1c�������i\1p/��pYʷ9���g\�9�g�s���ݻ@�B0!�n®�M�v��q���HHd�^.��E?�
1�tc)r�����7�$�7G�7Q#rf�)Ɣ�,Jj��Ƈ�d����'��`F�\���AЕqi|����64
��b���;������:��ׇ�c��t9�S����T����_�D�B­���FPAI�\v���z��d��D#�%������ <XlxVHYEB    3530     d40O�y!mp��eW����dJ��D��ɜ�g��94D�*��1�nUc�ػ��l}9B|QH-h������e�T��F�����6��^��\�pu�e����=�l��Y`t!�h�����H-����Y�Pp�ѕ�l��+!��F��t�7%L
��Z�_s�����y���O^Ā����4YmOE�T/)'mzLg��{�<>�K�����G���nL�_��t_c��P�x)�c������Y)V����n���V#�U��}����"Wl:J���	M�/�2��d�wi������:�J�-u[�ZYȵD�X�� ��hn�chZ.rp,��J��a� ��b=D��e�I-�!���t*��dP�OL�ݧ�/м��Jv��'�s[�����~;cO2r���/Cv�d^�.9�Go����9��i��#�~�m���pQZK�y��%�aw������~�$�Z��@U]��Q�����u8�ځ�|�]Lx%�`��~�۱��ߦ�Py�������xLPVs�(�p5��,u��T��A��r�'�8pA��Z���]m��,~{�~����%%�Qw��iUx���*Ѹ��>f��Wk�ywg�����Ri�Y/��ň���a��*��{@�_����ӈ�X�Ɨd�����NH,6��������X{��
]�m�װ�4���v�	��
`��lk���c��@��� �"#QK�n�a�U�N�|�,����*0\):/K�q���i�����3�`��Ap��5K{M����� �T=�8̀ɡ iU*����:N�����1�&'�#���y���l'[��P�7-}	�F��jN��[�fL�ϋ�U��[�]���%:&l���&c}ߦ���)��K���"���n=m�.RE8�}�E�*�,�䀹~H�9<�t�:C��?9��n!�"�~��q{A��G�޲��u(�2N��� 0sXR��Ȱ��C����yC�	���DU�LU:n�d����M#M�:HP3kf��[!"��굚G	�Uy쵓l���ܠ�����/��oy���1P^4~��]���?D���Hܯ<�:�vV�>�2�mv�ܚ}����\B�+8�Uڼ8�ȷ+�[S����ΆZ�6o���gF���\�����^>���!.Eޕ{�ED�b
<=���{ �<�O;������R�ad��mӅ��(��o��t�j�t��vzϿX���d5���@�ÕzЮ ��81�h�ȩ��5ܖ�X<��!)�Q�D��^��Z��e���w�S�]��$at�~z�G/�(R�Ӱ}�b��܏S�k
��������vO��hH��]��K}RĹ��~�����G���ݤ���'��[)�CG4��O�CYk��)dK�4&T�&޲Etu�ɐ���rU� I���n�6��L�4o����:{�/��&�;?�:�� ����w���>;�H��쀕�7�l+sg<�E���:M�Pn>��r
E-mz��ґ�,�50[��*׹�#NK]����w7��$��ɤ%�9<��k%Mވ��_d����Mds&�+B�]َӼ���᪅�����Xz��N�DҴ����g*m��D�|u��n���(�N�sm[�'QAG�>/-p����K�!w�H�-{x�9~��2g��)kbe��tÅ@h"�qQ��E]K�?��I����h��-d!?����&n���`��Х�[	M������o����9S��=���+-?A|�
q[����ި'�XG����'C�z�o,���`)���_�/� ��$n�J�W~�!t�%M7V#���ѿ��Y��*D*@���}�D,dY&X~�bˣ��A)ܣ�p�wd�-n��i�O�5a�@��cx���li[�9�������Y��:Dy"��L;]�9�Z���O��ݣm��KnA;�rҹ���+�R�.����6��� HW�|r�y�'I�5������+��K��l��<I���^�.l�:�'E�C+�ŎQa��l��R�Z#އ�/�N$�٭�-P*"?� ��A�xiz^)���C٢{�s�i��2�N'����zƯc�jӒ��u�Q~����:��y3���"r��l
�h7��bzW�c1(�O��g`�ew1�A�L���)X^�-�F�C]�/ �ź��9�>��w����u�w��x>��Q��!㽧(9j,�<6z�~:�~���1�s\�x�7����g��rdn�6��1=����7#�5��vx���d�w��,�,�
�ϻڿ�hX�v���65�"9�	a�a?�m��Ԫ���4��R��uL�����pX�>�0�V->�����,���B#����$Ɵ��=��~������~Y+���1�R����(�J�B�E�bg���XB��$e8PQ*��H/Q,R)yc��ݝ���Oո������x�֑�0*�AGw�-�Oh�0�-W؇0���k���-3�Y��k �3���#w�隍�3��2��dq�*�� %���d�>gi#}T����c�Ȏ��eV ���ƨ�r��?�D��QgW��#�P1��Tf��X���a�\�Z�/���o�����C܏my�����w*�p�/#��5-�j`���Y����D��]��u`ä*G�������-[K�?��}��Nw5�s�V]�{Cɴ��p�i��w�K�ќ]����t@�����]P���
A�9x4��i�H����U92�$6tۃ֧S/�p������%�������l*��JK?��wD��%P�N��'\{�[y���̔;���;�u�����b��k����1Xa�'�����a$T���H����E�υB�5+��G(�"ID���kH/�?��yAh� ���.�Z��Ἦ��|ȳ2-�a��	��3�kѪ�����`QgW���ɼ>���q�#�,҄h/-��	����H�ɕ���2aD�ⶥ��ǈs��G�	ڴ4��sT;/��`N������M��Gۊν]�헱�;�b���j��_��IoYܒC��.K_Ef��΂N����[LB;�����w~x��m��;ִ�=O4Q��-'�{^uT�bS�yO�hP���dx%ix~�+���ึ�p�ћ�Sc}2��� -
�҃Dh`�/��!AQ!.@�!iT��`�s�C���R����N��J�=�����忢@h��f9��6�����R�rG���\�	��I&�B�1?� �U�!�EŒj�X��2�ۄN<~�d��T:#m���

��f����Ve�����R��8O6�a�%�h�Q`!�j������[Q�Y?��j�$/�"����0�>zd���\!