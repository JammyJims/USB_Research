XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ʅS���]b�CP�/�w�q+���Yל@R���=������֍�o�=G�1N��!�]2*�E����A�G��p�ť�i�p0�}���#�'( �ɚ6H��0���1]:R ��I)�/x��.��KtmYy�f��Y�V��T�g�l}���K���@C��w�.�� ������!Kc�=";���6$O�o���X-�w�{�WXV�(*�����-^s���3G-ٲr�f'�I�3�l�_g���	t���#�pG#�5�N-c�����)���ov4;OV���l��ѹ"7 0�|���+{�fʻ�3; ��HXx���H[����KZu?�T�:nS��#0��`��xR���bc{xO��~��|�Ƌ4 C������d��H����6�.��(����]@���[p<��Y���B�YCT�H��dV.}�;;E<��h�<�MɌݪ��f�>]�߃����
Ch��!���N&����=�]����v�Ad���T�L��]�b^u��~�riݡ��xK�����Mj��.DМ|�|Q%/Q�����=[>��~#WR�9�ɵ"�v�dTގ��=�yM���x�u�:4�g�n�v�*H�b;����du�� (S�8_caW"��>,6�����!���s~#�������K��m�����W�cn�
�K�Ԁ�r�g��s�y=:�F�>3M�������=?yh�����F��
�}m�h}72Z);�<ƒ��N�2�MW�^!n"�4*��@�xhXlxVHYEB    2a5a     d70��yM�KŉLY�nҡ�F� 4��h�阑1�J����
;���^J�@�#�<�䀱w��q$����e��0���m�-^��~����d��QrlM������S_�L�/�d�����]��LOʤk�?�͘m�'�B){�J�k�h�ֲ�ks�"�Ͽ}�%X�Q}���X�F��*z~��F�{@��%�-���Y7�����U�fn2���K��Ȓ�s�X~T:��&����q�����6`�җ�����)(��(=΃{�K6�Y�>�t�N��%�jy���>�x��/L'd@��gX|��۹�MP�;��y��<#��z��u�Sg�?�v��̃�3���1�w�T��Ⱥ��N��u4]	w���ŉZ��>%��7�':�ZKzx��5���%��ߡ5���>��^��̵]��	 ���-�;��B߅�u���i%Ă�ʷn��tH3c�5���:c���-;FZ���o"�`�1k~�;RѨ��!�Ȑ%�z��r�h�q4�6E*�3:�à�G8�^ғl���h\��YYE;uO�.y,&����Z�g�]6��Q��il��C���~�K�H4��Û�}2⇞�?�<�nH}��s~:�#�A���_t��B�"IY�ˆ�h�Am�l��M�+VvVk���Z���#!Y��y���0�3��/�ɧ�ly.<7��#�Xj���4�iK��ĕK�/����i�Ie�eɢ����}S�^�;��X��{d����g��<dXV1��&��Y< /ͨt�RB�M�e!���k���+�X�&\q�g:ݧ�����.�Fg�~�0ލ�R��s�%Ʊ��l��˯Bpƣ��m���[AV˩_+b+-brV���aDtI�����n�Y����QL=[��A�D���J{�O8��bO�t*\��J~�s.�o�>�T��H�Nd�{��v�_�˼6Ā�k���m���|E�\�VN���q`&x
�q&���/AG�/ذ����O��ɷ�ߎw�O���Jgl��h�9�t�!�I��>EB/�^v-Ny���ӻ��<�% c�@��w&�7m��P���$�����h�_Ψ�t�#C�Y���r�9јzu�c�i�� "���t�gƷ������T�L��
zxA��.F_���U�I;�~Ͷ&�)�J������z�<�G5,�dzZ/*��HS6D̟����i����le�����^�i2u��^jKh����<���8��V��o�V_#c���A�-�-�}�<��rL��}N�A�X��kŦ���-��p���>���򕮡z}��9���^B=!s���7>=���~� ?�	�ʹ��ڈ�2��n�R�d&��Zb��\3��V��[�o*���#U�z�H?|�3+1��;�-!���َ�;_l:��ݡ��R��h�%��2 ^�oq����=�J�oRo{�>e����5�~�˨Gѱ0������!�$�)�ŻȞp_%g������uF��L8�R���Z����4��t��&c��iyC ;E���K=L�nE=������|;�'J�^Iż-����9���ѭ�LS���䲪xeEr�Ypa� 
I��6��R.<Kc�0#E����鐫Mݽ�<�]�?ZPDtN�5���Glzu�KH�!�-+�=��
�	�x��2�hc Wo��{kb/�q������O�\��O�P1-'ܷ݁RO[�lF����6�=�Z�v��H^J����A�
��~ɱ�(w9D�� �8�
����X�����P،�8Y�K��k���������͕3��������~^����'�+&j����ʩ���O���yN) � 7�ͼ��%eL�-��!��q@=mTv6�1�	�q�+J��Q�� �STC�RF�i�%}����_�}�'~�]c?k�$�@��-H�	��I�3x��:���u��=鴜|"_�,]r�'��6�V���ꑾ"]�`�־��H��nD�A���I�
a����h"���A>�C�]���c|)D@��[�����>�z�p�d�1�k6���"g�"g��a��ΌQ��*�f��o	��^*�iP1*5��L$P�!f�n��v��];CB��D���ff�`�n��M�d.� ͼ�t'�Y��e��� ư�J�5�AΦp���"a֮W���Y��K���l�1z*���g[��V��!ʋ�w{$�Ʃ��56���@����GMתl��*���L|��j�;�������ek����>�fUD�/���"Mi��D,��(���$�d�����/��15�lNEާj���IIX�6���?��*�1S�eQጆ���XrW�T����b>(����V�A�*�׶i4�ߺB
D�ȄC�g�Q����l?��q�'��I4f7 ��bv5c~�-�ǡ0w�l���x������?g#�/FΫ`Vd�^�-͸��s�mH�;4^c8����!��Dsi_�>D���A��;C���i҇�H���T��� ��T"�ծ��d����O�Vr�iw��u�r�F�a�?���+{��cp:�ԁ����7��Id;?�&G]���D������kQ%̉d�~���'b��,�K��T�'�`��,�[�4������9p�c?��yo7�G�zl��ShV_$�R�tb��W0����7��VM�,��g���ǭȊ��LQ���n&WۻO�$�\�Ϙ�L�Z��+c��c%{f,<�4��0D�V�ĈB?h��kb}0�ҧ���@��Y!��$�6b���j6B�wr�I��+R%Ca�1��mp榾�^.b������wB�N��Ʌ��{�je�<�����~�d�~�T5�;�B+m�- S��$7���x�1U�J�z�qMVܭ��Rb�=Jj���&lZ��|�q*�I8rP��ʞ��`�s�籿n�z^��y�Fwڢt�D����M5�%�{���=�V-*�4Q9�=.,�1S�������^�z�D�4*�gDF#G��.�f�Y��tI� ��z	�u�7�t��BQ�(��V��b9�Tg�
�QO������D�f_�R��H��Kc���ڼ��K1JS�ο�=���.-S����1�F�m�S)��4���e3��C�ͷ
sю�E߉A�-�U��,�_�c�6ˢ�_��Su#>I��HǤHIO��"QRB̼���7�m^.��u^�Ri����A�3��1��8���Z�'����6�����P���Z�/\�
b(N, @#���I��q@#oq��n@�N��ُǧ*����0��w�W�^V�K
5��b�`��]�/7�8�Бr4<���I��v�+m��\���~I��ށ�Hb�uAԓf���+�w���|�2�ߞ��腍O�}���Ds�*)�