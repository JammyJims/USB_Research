XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��aF�����}�1�8�,"^��Xv�A�Y+��-���\��^�o�������#��L6yG���: ):\<�����(�AA��䮸������B{;����S�u��$�u���/��p�鬠6ōOʉ�������^�I���<d�0�x/�,EQ��D��dz��i�]�|D*n}�y�����`-�IPJȒ�Y�N�Ă�m�`m�*}��LsbmWG���yؼ!nηS�]���,^�,_��jF|�Y�4�������H�"Ks`O,'�u 3vXt��EG7�/�JO�P����y��c!�7�Ï;�Y��}{=��� 咇 �����^��B�·���g�����E���3Ʀ�4LW�c��^��؀G/���{;{�N�������C�F��ɀ+�\�p-v��������$8�~>�J��z@�
���B~n:	��M��Fu�Wv6�h1d�fRy
zw*ڿ��
�h^}
��r?F3j^� �АUc:v(��)C��~1J��%t��-�T���P.����޸�L�R�mp��I�a�]�bֲ��Qo�&K��Mvh>������.�8� Ԩ�سX�� ۶�F[Xu�_�	�_�YM�����~mArG�@-=r\+�'�H��1��1��8�U��i<�n��R�0y%�O��y�ɵ��(�AO����{�z���ia+��)Dl���x�2~�J���>8�7`�yy+�^e�.��?�\XlxVHYEB    7cc8    11b0}Q?�0(�y�'������B�Xp����؉��g�	�sɛ#`s|�E�����P�E�� �=�V��9��i,�Ce{ةrX*���ɟ3L��!Ss��Wu��=U+S��'E,�Y�t6wwLd���ɔ	|��-w�7�A�w�-�K�>P�N�~�LRH��T�>&�4�(�|���;��" i"J��s�R�(n�ْ����'I�U�4��O�l��Ҥ\���EU���9)x`�K�� �=n#��Y�o?8����f����G.���:�d�y{�q��/�X�L�X%�T�KF��c炼�:$!�:�<�Z<V��+Å9���+����Y%������W9��;���蜮�=MWԲ�\	�����{G,��܍�ɎOA���euq��|�������ar�c�&��n��KN%D��n�/��$2�j#���kS��|�8��D��`T�; 鋃Ƿh�O=f4���t���˯#�-r� �7��s�7P��X\#/:���d�X��
��P�����$��[{*��v���
s�U��+v�VXi�~
����v�5��s���}5��y��ȍE&���ks�"�Nf6�e~�ڡm���T�c�>dRLsF ?L�`��/����'��%ok	˵��K��*θK��43��R`6�@x20�+��,	��2�M���5�!�\`<��4�mmn�r���ڡ��k����(5�<�qNh�������E�/�Gu��:�-�nI�����@z��Z�ά&�R����h�[:����I��\��Îy�du+d<3v�ק���(��K�������!\��wL(n����I�fAw4{%�=�[C��c1�WlqNec�7� ���{	�v6.�a�`�o�nD�4��;�W�] ��g׸U^�[����e�/��-<�*ŋ��P��H��N(�c�L3�s�D
�t�%�@8^C���6��j{�.��1��P�[ �t��rU�Gzr�e�,���^�H�>����dw�C�{�+�z��
�]��X=��j 芑HT$�|�7n����ŗy��ޥ�f��=f����$�$� K��L9��j��٬�UԀ�4hT�Q��0df��`� ��-0�%���^y�+
���^�-b��$���p����k��Ye�"���Z1��fBf�v�<�����s-Y{_��/W/A��=9�Q�""�!qU�ǐ�b�]�n~ն!B��P�M>�e�J���GXS�I<h�Zaċ��L���ހd4.=��e �e�2�\��_�����H�ѩ�SN��Y�k�O����b��mW3൧��\߁=�����rQ�H��0 �b�~îi��5u��-��u�.�zb�D�7��zg�q~�j~[?9�\��2G���e�LքA�A�L"6
00/D2Z;+.qV>y��	pku�j��c��s��c�����%������TY������PbO�����~o���<�R�Z�
_u*ZL�>�v��}�x$`ZJ�9)-\������-�<�S��.Aa����\��+A��1��V���L>��0�#���ؽ-�]}I*aT��=��S���av����U��f��L��V�hgZ����V.IQ|JQ�]��21
p3�"��L�|:c{��)�HDՇ�!8��d/���Z�*Ef�qbN�����;s�Bq`��.[xB��pF�O�M�$٧TҶȥ���|�q���o��{؛g��>tS�v v�D֒�L�0u)]���~w&t8<󜏙~k�S(��m�2��f��n$�v�&��&CePӑ�,Q�ښ�a"z��T�P�����X���4��%�T[�7���8\lms��R
��A8��|�b�j�DIl�K�y܉�)�<'�:dxܚr�Sxt�G@�k[��+�jP����6�mmD�j�^�@������I�R�K���\����Z��Ȑ��r�`�yf(�^ʧ��,�q���h�mf� pNȶj��k�����.���Co(�d�Y����%|�`��f��$��;���y{�q�K
��ZQa#���>L�����~o�28���=_�zj�Z���O+~�rB�W8�qȵne@��ǭ�H�̲��z���C��쾝�3H�ՃZ���7��h֮�h5(�M6�]�O/���%�ڵ�-�+��]��/ZT37�0N?��5j���]��A���\|�*�L�_��k��撎1ᬄ��h�|��9H!�iZ0� ��&�ˀ�uϙ�N܋N
[.*�s��H
��3\0Dȷ������̊(�t�14*��6z�*i�N��9��mΝ�%�m�T���x�ȡ�Pv�Q�jWP��ͬ,Ϟ�0+l�{��qoH��������#��U)yR��i�js��p�D]MJz0+ԁ�l���~���̠��ח��d�%eZG8����?��A`ǻغ�~�JI�4��q ��L" ��;�b:˃ֆZ�!���Qk��m��^O�{$�̹
���8E�m[A�pac��e��P�@ 7��!����;F��q�㳙�ώ��G����eaڀ��&�����
�;��:�.�N�i|*�t������?��|����[�!db��i��_��
�9�^#aPcϨ�cN����c�VF�:��<*�Bu����Į�H�����?�a�����1a������z��ߴ�U�����������yL|� �_�;jϜ`�'q��L�I�l;/�b���Lj��0ϙ�ow�K�>����k�����X�Y��EJ�uA�U3�jVRm[�N�*��ڇ':���]�mlֿ�ˬ� ��G�֕:<t*�O�ˑ���� ��2�#�(�^�r�#U����ƒ�����W������P?�b�R���}E��4��܀�П���<.r֞�H�w�z�Եg:
a�Ղ5����qZ��ɕ(��aC��S������\���ߙ������>����r�z�g��lx���Y�qgm�?@�9��B��+�O�nб؍<
)��g��Z���1����H�E���e	�+܌�M|���d��^��]��L��� 4�QB�m>����@��Lvſ��I�/�`&�߾6w����H/�������~�4�l�,�����_��`Aj��Dx�`rL*��5��l�
���av�l���>s�ˎxŶ�ꐻ8� /c8�:�g%�C�I�mw���E�s[�V)���W}���c2���وI�K} )�Qڛ���G��-���&Ʋ�.���R���QXv��V��#WC_N�J��)��a�Q�/�J���͞��$�vl��X�Uʚ'�Ҷ2Y�r,_̖^�r�d�:_Wн�3ۨGLi���k�e�r M���O���RĖ����2wxGZ�:sO������i�$�Ռ���R3o��t���R5�Bg�iC'������rM���`�������Њk����Z&�N0��zr*�a�6߭q���	~��-|;k�4m����)�u���m�����'�?�X0<^���2�x��iWs�����E���ˋ�E�\V�s��:�kSϪ�4���F�� ��T����/�.2i2m���S��������A��S̓��uސv�P�$���#�X��n��H�HƸ�r�V[��6Y��t�V���@� �L�³`�xy	+�]9m�HG%oY��T�r���]�9"y _�^��.�Y^�1�=N`7�|�S���Kl�n����w3��>D�o�nL	����(��"�D�~L�	�dZ�M��gK S2Z�j����1�3�V�����i�y�d���*��h] �������1����H��];��@P�q��(��R	����P��C��M�)1�6�̊X⟚���ԞW�LN(4ݑ<7��.#T4�|lP!��թ9��E㎎�V�G�R�����Z��	���+�n�-��Hn|�Me�w�KQ�M�oLN|���#U����aW8��)�J����@�$J��C�����@9�g\מ�?Nw-+�#�����>rx�Ǚ���bnS	�U��,���"bgo�ݽ��!{�H�-�C�p��Y2�\�/�@�q��Y��Y�2����AI�>7Q9����I�r�y�@�F�Ĝ�-1��B�h�����O!��A�Y�O�o��LoO�\�y
��:S��(��%�3��%B���Md���X7c�+�]Q��p�Ǟ�yG��������"��U���ґh<��s��F�N3u��Jo���Mxֶ�8�W�$����c��,���q�U��FF��������u�u�Pf��,�;$�ov�Vfb��GXV)�:�
j0if��@���>?�����Bs�9J&
�Rr��)W��dRw;�Q�4�|��$���C�`\��BNj���-�n��[�Ă�zx����駡��Ĵk3 O�v�(�)j�Z~\�����5v;�}�<�eˬXi�{U]o�ګƣ��Ar ��F;*�e���$�j�'a,�Z�
^'����gL�'�v�B��