XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��є�Sm�Z	��9�$I����BiA���GY�@�!G����Z������k�y�$»������1N~�� 0�c2�j2X�@�����T��@|u�Ҝ�� '�6��e���,�_���ǹ��01�(͆�Δ��.�~���a3(h��;�ƍLvl��A%'�� H.dSPs��6�X
rҖ�j�{���5P?�C)엙%Q����O�;R��z�Ht�Z'��F���#�=yh���#7��,�����Wں�B�h�"�rpJ{��Wt`#�1B����E3���f���ZHO�,�r�]�Y�w9�c)���`C���;�"nb��G64Gy��1��[�I~���$�Z���@9�禣M����M2�T�T�q���5"kF��hJ����z�7ꦧėVթY
�h���,Y>p�ĭ��E��9�Nu��#Ul{����,v��/y�Mo1ɃR�w}ȻJ-��6�b�	�|lXX̅����x�����t���Z�g6Ω3<�������_&:J�$F2�'�t��(�f9���IJ%��OD�x���JD���X�)�[�B�h���)åe�<��0?�����q��tþw��� ��j�`�\f�7(��>�����gTu5��y�8���F#h��s�>%M�lr�h~�pE���M��+�C�Ð���LB������.��Ƿ��Fu���o)��+&����a�-��KB⹱��Mo�M���i�^�0���G04ZwP��|2]�}��rAɿ���XlxVHYEB    357f    1110�]����}�]����(�8 �4G�@n*�1�ד��y �L���8��Z�>pp��8N#�V�H5�%�����wB���p�X�e��Y~��h;�����z��4���.�A��E�ᙃ�Z��)8����JB"�'��u������&�=mI-&�E�ML]��Z����l��'ɕd��Çi������"\E��@p�6w$����B�Ce�	O��ErNo�������B�ccc^�@�gU�s�-M�����i�����̐M �ȓ��u'{߸�tI	tt�1sǝtsa7]���I��Z���E�Av!K��Ar�^V�=p����E"������Q��jN�d�!���$xjGHXD��Mu�w��s�WSj5����������YFrOvP�5^���0N�6 �ky�ҟtn�Ya��D��&1g�]%8��m5�a��r�������n˲.��[��`rc/�t�+�h5D7�C|V�@F�CSa�E�:���Og?N��82�zV�j��4Jו���p(�T��B��t�5�| 頎���c?Z6`$d9A����Uu&���fw@u�3;�{+���tJ����e��/Bo�aB���Av��O!�� Y�]��N�#c�ނ_��Ko�D��`�됇Ǜ��	��U�)��
K�Y]�f�\7_&x.�����n%�;z6�%���&cߴ��b=�Ϣ����`Ycj���Թs]v����I`���3��������M��)�[�c���1t�\�K������:�?��3u�L)zJ>c72(���OC���hm|�nO=����iR��dv���T�~p�K�U�^@�L��>�dxP~8��0����4��S0���H5��.�<gCv��հ+(pN���p�b}/�%��_��k@ʍZ;��Ж�.�����%��F�-F�-��Mů�~�_���蔩4�}���+��.׈�\��ҡ^v�mZ*o�"��/��S�S��.h�D�5:n�,$'��jmh�tƅ���i'Q��iM.�M�4� �h����x-+�Wxu�~B��"���i��x�i��9� ���:��W�d,s�X�VF�ddgk����ʱ��GN��\ڝ���4�}���D���/9A�تF�H]��?�C���Dǯ7�� A�sR�}�����me�F�����ώ�o�\=XL5���^o�B��hq�����ܶy ����J4ĀX��V5��g4���?��%j�'�}dڒ��fLb;Ys�Ly�ݢ��;��(�}(��R�F�!i�,P�������u���+��5��̗�,��v��=@���h�m�Io�-����v�[�y(��꠬�^����~�a�H��*5��X�����s,C|xHM^���+�+E>~'�3,�< 5��_�����_8ڣb
�-5G,���=��B��8M�m T�3����uD���� 0�:�ΟN�7f%�!Q\[x�����G4V�sr�]��{��?hT�8����t8n/��[B؁y��	�nG��/ɰ���*�p��l~�Pb@�Bu�'b����+�sF��H�ȳB�xHZe��\A�y8�+~�h�B-�
�����V�1���ā�	gmq'�-�b3��B	�#��іf)Uu��ȕ�	�%�D�߀@�VjC4l7w�1-+��]eE�7z@��2ԇ�cI��	�x�8y`�C�z��=��!Ls�<��f�}Mƈ���{�JP��������O��ٿ{����Xr��LS/����Vt�6�r 檸���D�{n�z����Kq�I�������� ��^�^T�5��Ӱ~;A�ڄK�l�Η�>��?��j�b�u=�b�"?(K�C��H���l8���f����Y7�l�˺�ץ�ð��������q���z����;��a�?�q'�[�l$��Ŭ���^�PK|ryƳ�/�A�݋�vfa�G����^��)�t�?O?���������3��Q�۫�N��T��oV��DdM�d.��� ���D5��`�(FO�b����$�"ej8x}*{�2dIK����z}Y���MRn���Y�ȫ��ǲ<�<���rg�ɺUY'Щ�,�\����۵/�?�ȓ���łM����+I�gU�
I�i-@ȭ�̉jI#q�弿)��nݬ�����+��"x6�qrm�i�j�]o����\KP���N�g_��sY�c��*�:`=⡣�D<Tx��o���Bo�����>���Ț>b�ǹ���4�rP]L[VLTθ�?$��Ltͣss�J	)О�q+	�=��pe`E��i)��D9�UAd_l�*�������j��5�ڥ60$|�5s��|U�������az��rF'EUH?FE ̂eU�8#M�����Y��}���n����B �N���#���g���@�K9|�Qc��3=ק3��&��t���`��葷�i����bjrrΧ�����1z�D�	߯�yl3$��Y�59�F�rFK��+���_v�P����8H?�݂[��*�S�`b�s��a��HxYzHm��"���}�=W�vi�6�̹�@�AZ�7�����{�!��W:ZJ�ۻ�����a����dIis�E��J����˪}s�!Z2ΏN�T'wg�#K�����iu��~����!�y��� ����U��O��ey<��Z��9f�(�'T��2sE7��'���'QBZ5����j���6��x-���Yp
����y�U&R���kUTM# ]��h֭xZ&��� �W�}�y��&É�. �.���|���DOE���3��cP.����8N"�F����#�S�UP����ng�s��8�9S��o)r��=V!�I�����q�4|���N6Ƚ-K��-x��Οfφ^c�5������1�*}�B�7��^�:��s�y/�d���!�p�.zԦ_���闁���i��>3�O��J�0��́~_/W+y�l����M��-e�Ûa���j>�Ĳ-�Xm}�H"}�C�l�K2μ�܌��˖k����zYv5(G�F�}d��ި-��U�.�au�55à�`�w�h��9����M��Ej!j%�u#r	�8�j���e��s]U��XbS��a{{�D�,��9|�<�
]�u��z؆��C߭�x���=�kS�q�0�Pf�c�r�@�
>�"��Z���am��=kpɞM,��{Xw�F�3�^�3C3��)]|@�m���)3�!L����Z:�'
݆��l�~EzWb�ujo�Dλ���/-ɀ�7ƌ����E���g�徝����2�,��]��w�9�F>"��郋�x:	tW�a������;���\G��O�AO��������Z�J��{��:�)�Z�=cֽ�Zs��	����a��4k�L'����lwX��Y��.x����)q�hq�m�V �э�܈�"O�(��^�z�lP"V$�n!���DH. ���?/ϯCc[di�gi[�GlZ�@�3���C� _HW��p�p��UJ`!�d;�G% _yé��
��T�
�)����~��=�FP��qUS�}^�b$p���`9����j.t�������3Hʞ
!8��!P���R)*�������"�	���{�(#h��C���U��R��������Օ�F�]%7�ړ���w²�+&w1�a(��d!f��u�
2�!𽇴mzlg^lH�ѿ�T�]֜��\�U��$�8�^����V�OK��[غ��"�>�jk��|��Ytٟ	��%��i�6���I�^]��|Mѯͱ C���_��'�j��!���-9���X��JD�|�Vd�ʵA��a�Z�{Qǧt83�S��L�\�+ �b�L�e��d ���]�B�D�d��/����(͕[j��h����9/��;۳��pW��O��^�Hᗥ��`��U`�m��ŗ+>%���8�c������B�Qd댞�Ֆ��0�2"�.Cσ�
r [��4�q.�v~K���&���{s#��A���Ē7�$�Fy��Z��ȼCy����MŌ[@��Ӡd�Eʖ���	)���F�9:�0~-�?I�l��(y<5����%*}�N�%��u��U���?���7C���>S'�dz����pңz����k�"�:~�+�
��|�\�7'5=#�@x�\�ض��R#O��Nb[�Y���6v�$SGd%8%}��B�W�&�=Ov���Y8q�k��;���W9��#�P'On�z�jR����X	����-G�9�