XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����}��)٣�^��օ��r�T�}�w�@�['�/�d&��˷mև�z݃�L-�!z+~ʖ��o.����%�3��x�Ч_��PX���#�"x��5 ����@��g��]=c�,�H��J�Xm���\ʡ�C�!qlV��w��&�Qv)��䓲~�<'k�@S�~yg=���qY�8Z��X�RD6�}k� �	��2�5�S��׷x��mN�Sፍ�D�J���,�`�r����� �����؝g�-D�� 	b��˥���+J���c��L�>S�h�d|���
�6R��ڣ��c����	i����KI+���*�j���7��p����#�@n�@�e�d��.�{�y�(��`�g�ԭ����7��+�[]`�?c)����z�]|�@���2&�D!�pϐ���_,�#�̩��@pXx	��H��)AnN�%b��hP4f+r �;�o�]b>ڷ�\�ƛ���Ж��~����Ã����h�i�(Bퟮ�fb�d��O7J��2�m���f�l��|%��H���d��+�Y) �Gɰ��4)@�6��z'�p�-�#3�h![<�Y�1P?l������D�u]����撫�/&D�Q�����K)4�0G��!` p<&̥øm�������nzP�o��D��g�/Ka�c�ƺ,fh�ʆM�y�i���͵_��?��,KR��6�1Ŷ��ڞ�RJ3
HER�Pi<��-�Y�����~�]���[)��/r-�PC�|K���|XlxVHYEB    b2b0    1b30ND �j3/	q8�͈Q2���.�q��	BV�r�G���72�z�O}b��
��� ��@�� �ؙ��e~V�g�(�9Hb��n.'Ic�:!��3��2�Cc=�3�胾�.8��͹Ui�i�B�'��<@�rq���슙�)���k�<'N���ٶ�h��j�!D,�+��UCb<��G�l��[mI�VIk�\�(uE?t6"C-N1,`�I�o��a���S��O�X7k�����"����o�<gm��d3b�d\��e����KM�MYaG�f2�Z׌5:�����)�6.��w�����f=�XR��@d��Jf�$PDuî"��[��U�h �����}ýO�X������E(���7�|��q�� S�O6�����P�b�st2=�Y��ml�iK�rg��i����en����4r/�JפƤ�T��u�+��I�����L�r�S�S��T�P�"�
⌔��P4�=qXu�l��9�K��N��Wr�đ��v�46�����Ђͪ&��9H�p��V�:ZN�n���W=v�G���(0�8e��F.�����TM�!�2�yB��`{f"Ef+����,^��ݗ+V���I�a�Q��`��K6_?")�B?�E���E[�L��7�G����� wwB�k:����6��RO���4<�G}63σzLT5�L��G;��(�X�W�fb�ނ�b��{	���|�A)�<g~u��#>(N��p?�Z�_��5�6(���7�l�/�s �Fع5�עƊ�#<���1H	�dw��*1M�Y�|u5-{���k���~= ��ަ|r����Y�<�CnEː��U�#���������v&�?��N�%ʞ+�<�zMb�[[�C>(�f�J
��L}g^�	�i�ˍX&�v $�a[?I�$:g��2)sn$4��)J��5d��iti��jE�r�>O��u�`x*|a ��Ű=	�i�_)M�����f�q���=ۖA�f����;?>hO7���$:(Y�K��'^f�qa^��a����ɉ}S_�e����N�<�;N�"�+�2&r�(���YhS�ʉ�1F>�)���N�|<�׎hͮ�c�u�~�#E�g�/���Ug�P��M��,)X� Ԧo�K���( h�t^;vN�[�F��{��L���žv�54KaV�
�^ "*գ-%W���[��S�»�te��@��T*�=���{�jr���JS�+{�������2�&L`u�Yjg�����\�@(��/N�����oRbX�cY_{�Cr���d��țݦұq@g���46C�o�BuW���7 ���wY�YY>�ֈ��%A�Z�5����C��o�M�*Φb���߯���g�\rƭC�5���}R�Ͷ)�bV�xi!$N��7T�	.�TV�%-���O��[{��!z$ů�ߔ��bBD,���;>�h(�Q���x��V��|������Y�3ʨ/�&��-�S-s�E� �����H������v��\_mYE"2��sXa�{.�<%�JN&xK�+�6��CWKY���H8k7���Z!��A����~"	�Y=��zȁ�O~0���N�\�R굱Ϥ�t���{��^���uk��N}C�t??�3�l?�k&�䠉8�vLG�>���U��L�߭ni'VNe��eH�#�"��>[�57�Brcg�e_�	Q��=�-4'�����0�����U�N�D��!��mѥm�����|�f�s�>;h���Κ�(�R.�6�3�M�^҆�!��'�o��Iq�����%CR:���P���g��C;f|�
>��G&Z�y�pأ�ڝ,��(�f�݆��6�LR�I��·�W�c�m�6g��27ו���n��#).��1������J1��y!󠲅��R�cj�#c��`C@3m��'�C���+��
��O�;����Nai�q�=�s;���3	�%�]:���!�y�������,����_X�B��[ {���(g��Ό(��^��^���Hi��.:�эS��(x�uƬ�|�m�b��������O��s���<�9~ւ�L>j����$	���X�*�B}Z�
�#�S�q�D��6��{��&��k��ЀcE��xI���g6.�d�w�_:�lg���P�a�:�3m ��W���$��%p�Ӟ��L:7�	[�0FU�����.�K��\�Z��׊�Ɨ�x��b�Y�YV�ǰm$����ȍ#m�𸉽܃�߸�'+�m?��ޡȸ����NWf��CMBӫgjH��V��Wǲ�I��KD��|��c���`r�nx��;~�Y�-C��(�� �v�᮰VX=C(<2�V�~a�l*=�6�`W��C"�1�n�M���p���g��0i7z�'�r�'B`|����k4��2�^�m�6�*4p4J6c�ަ�0o��I_�p �5�{�9��ޖ��8�"Ѝ�L�ߔ >)�Ymd�m�u�C;��^�xI��KC�g�����m�(� 9B�3YHP������z��lf���\ܱ���!�)�jT�`O>�)VyL#!ؿ| %�M�A���₾�to��<��6���cxǣ�7��yϘ�$���� �����>ƫ\�z�8=���/#\V ��	��-��.�n��%2�/5��}�*,��)�"�3�,jс��l9C�v��xC��wKl����Fe�5����ü�#>L��a��l
.A�=s���Q����w�-&|c�VYT�v�x>�d.����<~S����>i���6�Z�����2qu0ĥ��q��TA6c�(<aU9� ��&���F7�6����A�i��ؾ�J��*�+�*����E��h�A0 T�09Ij	�GUȓG{p1�<�;����D��Ұ���g��[��-c�������Ù���]W�y���5~�����l�S:�A������Ap,�� ������0��-#�H�Э��! h�EzY�2*<0.1�Gn��0���d����0��/-:A9�B\�Y\f�6��!_`������ٶ�V@Njw�U�O
m�
E���/ht�u,kyҼ$ٯ$7�u��A%?W}�{�oA��?�>]�I�@}�����nys:�\�rՃoc�Mͣhv�g�.����^�K�����y��:�jp����Jj�������B����L�g���1��˗�C��i���UWc��|ȋ&kǗ���q-7�y�=:��J���Mj��-�j5��L��I�_d�_�z�eh��.�'�.�Pgj�k�BN�#t�N]P���k��Ń�V��6��Dr�+'����mY��ۺ���F �D���U����b\�����Dǚ7e�Rx�8ų�3��gM��o�TaA��Ѕ.%���Cn�W���Ӕ��_!�(X�|׃����QfU���-~��@��iƺ���G�ȡ�� Y�>��M�fE$��m�Ї�/���l�k�kcC����Z�����*}��W�D��ɴumf��GZ��}C�Y)L0������Cd3�K~y�k��lZ�������\��+Gy <
/����q�e�tZv¾ ����U��6�:�l��šgv�3�L+�K�U�
A �Ø� r%RA׶E�6g�I4��d��8U�67J ̐j�ɡ���6<��p>l .�����"-�*z[���"Ŕ� o-T�m�X�Bʏ
5�5$m`Y�uiT�����H`������K��^~���"َ}�+�g�i���#�g�a��u��!��;+�Ї=��Y���Jt�Y��3|sLfs�BJ�xfy�ӑ�^.L~#wz�%�Q������q��J<)���X������$1�����$����ܜ��"��{H����9+�ŭ<����T�`ψ���q, ��FLEk�]�y������F����\z���*���ڦ;���K��	�j�7n��Juz\)^j�#��C$G�'�(�mA�����2|1[�Гޒ�`F&jHt��7�r�D�E�鱖�|�����52�f �pW�%+�}M�VJ�)0T�!�o�@�_+Ol��0�q���Jw��7
��l�o��z.5�=�/I/aC���pW����Y��K���*&65���tz �i�����oAB�z�b�1rfn%/m��=��i	��x�+���d4Z�.~H7���� ��U����F'6f�bU�A�z�fT<��B �[8h*�Yz�I��w�6�u�0������?�M�
�� �A��l>$8W�����If����?'ЛN��XA��m�8���Z���o��y7�i?��Gi舟� �!����o�x�宐��߮M��J:���Η�B~�U����T#�4mP,���0����h �`�R^bC�b�1#>�/���G�$ �����˵��thVss��Z���gܪ����W%gr�ր��-	�S���i4�S�X��t�i0�-�.�*�T��y��R?��^cS�n��>0r��b�d�i�[I�P�S����R��>7��m��( />�3�J2�P�,���$�1'ٯ�+�Y��b�f=FI�?)�|DB
��OI���p1'׽��&&c��$Ot�摵��` ���F w�u��c�̸Aٹ��J	�x�#f��@����'?�����|�{��Ҡ!,"%�eQ_ [&��Wx ]�%�U	^�,=��G?f,��`���h`��do��@�f.�<UCn�ߓT��԰�矞�.g��Yc:�"{ ��Fd��U���YH����'���v{��G����P�c������X{�� �`J7�
�]���`T̪C��ac�����	��"�q�y��ǰz��N)u��������6��]!�=��X���l^2�5��rȏX�#�w�����v�Cg�O�$�'K�Uo��]؝X��;�+u��J6�V�N��p̬ {6$if���_ξs��}���tl*畺��m������t�9L��W:e�a
��U����C�܃7�b֛�B}�9�!s�bK_')�@eY<��O��_U����r�U;�(m*^��}4�_%�E�5L=\y=M��>^�q��=f�-��.MҦ*)Ǉc�w�J�D�JH���(������V�K���z�G��4��%�1	�3_bn�Y��J<r�@F�0{�͜=�Fq.h�/jW,��´y�1�sm�=���4.d.~��1��F�.�a)BNҰ���w�,L�AF���*t����_�mf����	�&��5>��A&��܈Vs��a9}�����IT�w/�6���d�Q?MW}��"G�hr�x��O I%�	G'a*^��+pƦFFĮ�Jěl+�����0��;���;�ȸ��E�HS4����9K ��9�(�-&P��^��T,qȹXŌ��*C��.!.��@%��* ��ݮ�ƀ���t8��n��-����)L�{�Y1��e"��E �y��1Bc7�d.k �Tv��&O�y�O�_�Yc'��+%^�[-�3�\���N|��>�OU�p����go<w��R���-j��{��8L�j'��D����/�?>���q���yВo���i(�Ű.A�\�Q����a2A
talg�d�J�}+��W�za�+����qY����bh���Y�-���ŝ��h��E	u3�O�a�(J�OB����4������su��K�����N���ϔ#�[�a'F�k��2�3�B���������;����S=�ᨈ�/��|��M�C�7�Y���ˤl��!o��|["��gWI��A��2�T4Kw��6�mh���GLpI�&��4�ү�:�O�_�]�ґ;�P�D�k7�V�d���Q���C�F��噙���5���G;��k��\�D\�$ԕ٥7�˿ihrf�k��b[M#z���) \�:��=�����"�d~�W�顂������vN��;��W�M���������Ui�����Z} Аi;�A$��VQQ)��[Z���
)[	1£&�b�u���F�H��D �p7�e���۳�M�M�����"��<�D4G��IƮR��\�Je��D(���ѰD<��+	�4M�֍g���[�:�䜠)�b�T66A�N;�;�ɖ^�$��1���p�˝s� !�h��_)��R��K)�U!�����Α0Z��l�\/F�Jͫ���v����Ϝ&ZYR�tR�}g��1\����j����,R|m���R-,�R*�#�O����*)��g��L���Y#��6}N+��"	��T� ,6VB�>�.$9 ?~�$
����˳�n�R�����(�V���v��X��9ܛ8M�mb�C8%V�F�0�-*w$<G��*�3��%E,+���:�9z�
��OW��Sn3L J��&�O�=	;ˮ�2K�%�6�U�&2W�f��mC�d1a_~(Uq��A݂fiv��AD'(P��T�z�Qү]d��1~4�Ap��Zƺz�H5xdʍ�J�Tf���@�AX��l�*�~����蘂������d$��<�=*��}97�[�	֤XY0��W�j���m���7�gJ �PUA��F�����8��l����׈�L�_�M�@��#���4(*�m��#���]9T
�7���I_@X�J��{i/xFqu�����ۡ��04Y�,��5ɲQ����jfW�oDIE�\�b�np%,>�v��<�_�j����E8~Z�'aL�:�F10��mp��|/������U)괍���_�t�-e�2+D��e]��������xh1�92|t��{�o�i��~*~
�u�/���5u"�U���UX f%�Fp������e1�
-m