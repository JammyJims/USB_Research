XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o`o($(�1������*�w�&��$�l�ͦ�1l�3qC���zA�b��!����z鐵�! �I3:G��n�f��Wzw-+W�H'k�W�K�ө�B���<�M@@x�5����8f*I�9�w �RDK�g�y&C�o!�å�L3��	(',�̲�c��K"��Ч��S��^�;�c�^(�qT����]��}eې?��-$� 4l��籁͎ �uW�IRP0J]vg.n"���f�.<Q������3�����<����%�mb����g�8�Fc�͈��h!S˹�7�0�ʔR5/�xr08��zG3|�2�(b^}����u(G��t�ۺ��N�B3�֤EV���j�iy����\Q&�hTǄ�DR���f�`j=*3{�r�%?M���'�\���	��ݟ�o���B��X���0	b�_&{=j�&S�}�)��5Z&� ���Z���`@�He(��],diԵ�hTf-��I��B]��O
���F'��`�@G"xzUdh[��G��%�9ʥ'w�l*-L�Ϧ���B��}���(
"7�G��!�1���-����b�#��r_ɘJ�����P��a�C���!� b��2�VD:D��q� � �vڜ�Tz��ד\x\5Mk^sا8H�ۛ1�q ��/,���}�����̣y���o�<����a��ZA~=�WM]r{!�(��HH��e��ۛ��j�h�BB+٤�־���H����~^<@d�՚��XlxVHYEB    17f3     8c0��x�C�䭽o��NJ6����q9�fw2ޕ��!@��c��������@|���ʷ|�AףYɄ8n���G�dmy���u��r�g](�Яep /�{'�/�:���y�44�)�~a�׀9��9���x��n1j�˓����@b�U�]�`��X�v�WX.=�!|��K�������Q��*�Vb����'w�J�l"�t���*V�5dnU�"�"�Y��4�R��⛡>D�Fڍ仰��`2�n��ЬلjH'�%���
��ب��Ե�@b�S��!~����R��i��!b��ع�ӑ��˄���-93z(̠L�j��锓AD�˒������j�˯��w��N�`V�B��d_ˋ��o�q
o�"�\���-�S�ߥZ	��~7��i�r7I�wxsc��+�����Ǯ_tT^���Ys�A���,�����T0n@�l������O������:�@g��$�w�e2��9��㌃�3��V���7A�G�Q�1Ba��WXH@�.��toUk3�?�j��Rg�3ʋl��r�x�����_O91ء�?�܊A�
 #QF���G@��?�{O��1m^�9�s�/
"Y���K�YfA�9�ݚ�n����������r���r�og���ͣ�1zO ����E?U�mu	[�-�Z�?���3�T�ckD�髄^;R��<������tL~1�;YH�����d���i�f��zAe�iƪ8�5�0" 7_`*+�T���$��4G3L�AuV�'0��BDo1���//6�{�6�h옞�C9V®$�JЭ�����PE�C�K�a[�P��n����Z�3��~	���d���J9��؁�o;��k�s�W&=w�uQq�ID�ծCmw##�r��WDe�#��$�6P���]�y-���Z��3 :�zT#�����5ns4ex����-����h�Q�8��鏗��A�v3�Ѫ�hv��	c�49��pr	G%�CTFVlWγ�@�N[Ί����13b�a7pQ���U�W|��uY��U��k���8�<�y(	UL���h��ɴGK�I�*�Y�"����LVy׉�w�w|k ��Q���3��#���S�������%��v*������Rޅ���9�g!�@����p��aΕ�^���b�3���@��N���qՙ��;��l�V�qȊ��c�$�p�6���/���U"�G����cD>^}� ;����`��J3n�vt�`y2�Ҋ�kuA��lCCIj����!UKӡ�5�Ob�x���7��,��T�Nk�xd�:�O�v�]�����)�7G�=��{C$�>�0����]Q�����Xa1��zY��Nܦ�������q�a�R%3m� ��;��ȃ@w�}]��x2sb�[���d�4k ��㸛d�uw̾�S9���}�Z��/�C,�g`	fRN��	��=E��aԅu����c�Kb����sڝ���䪔6���f��*4�'�#�)T�UI�^؄p�.����7+;�sjχ�ш䋑���%�$c��gr%@Y�ߓV}Ѧw���#D&b�n��W���4+���b$0���C�.�����{�,�X�\!U�G����⽚7�g�a�ȫ��Z��z�d�@:�*����2*Ȍ������(q��b*f�^_�d�%ݣ�e�8��a��Q�g�B%�	��Ԣ�����>L=��+����%v��Xc��
��7�ﺚ�M�:(?l�����ʔvz�έ����Y� 6kqJ��Q���n��lZX�Җ_qʉܪ}4�7y/��L3��Z$�͓7���g~�+�'uӌqEX6�PV��ZJvF4U�(����n�05Q�-��\B�|~� .8����o5{I��쥽�L��yx�&��C+8p���	"�)xv@Y\������bB�-QؘEò�{�
"���s�2*V!d�y]|Ϸ$���K�[���!��dM]p�$���
�Ttw��C�2S��x���x�S=)�Uɟï�5z�Vp�$�FC�ר*�b$onz��3W+�˙`a�"�'��&f�L>CL^%�O�7o��Ī!]C�?CHr�$2���!�UHF K��q4.q�z:�yr��p�+H�p�J\����&�K��%D1��C�gND� �iX>�È�z�^�gA�ty�Z�����F���q��K̤%Z�%,