XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,����n�I��%��2F���t��~v��`��[�]L�z�.7�wޝ�*��J$�̀�d���TN0�� x8(�J���+�s��o�	�L�Uyg*��80�����3N���|y,Ꟗ�����w��쮇��ͽ�J��1<zX�y�l笪�K=$�6���nO*��9�5G����p�������'��3� ����!9dSHa��l~�0LG��C�K׮Y3-�����P9?>�f	9��z�=�MS
hx)�@��xr��s�'�KN������-���e����U��vY/�O�5��7��ѰӇ{$�,�{$��a4a+�2��?��n�Ғ�@c!��ܷj�S�����4OƲ�d��%���5�H�>�.v��7����L68!@���`�_fN��}���ӳ��wM��3�w+�BY)f�E^�*�g^i&��M79������Ҝ�A�Cz���X��Z]�x����^M��o������3��n�@�1+I����\�Ԣ1{{�:)��Zm~UU�}|�����ल�w�ۜ�%��&|��W�{�v����:j�@�{̗�̖��Y�T�."�����Ñw?��n�������&W�naM�e�>��_l�I����n� ����'cI={���M
��C���F�_�6ﳶ9�sY��:4IGa�hM�/���mE�����r �>�HI�^�T�u��0�B�����!��j7Q�(7�՘��e/��6�D�'������(#9�n�����o�XlxVHYEB    7ae9    1aa0�)��5�ؗ��.=�z�"���{[rV�SW��E���e/�}�\gfE�7ז[-�'��۝� ����ƚ&Ţ��&����HC�j�z0�=ꎿ�/x�}Cִy:7��(� ��'$�ZrD��A^U�؀a0A�k����Fgk4��8 �)~	OV��Wh2���W�C}�����I�#k3W��V�	H��hٮ�Y4�zD���e��W�`!�DPB�H����4�1��b�H�$F�"Pc7�B�&��>(�g��ǎ�[�+��D�h��s	���]�f�<��sYC����'F�����| W��ߚ"w`���ÏL�W���Twa �s� J�2�c��Kf"��(��1�v�Asl�������^i�:�3(�+y4՝�ΊG�E��Ѱ��R����nA�Q�ث��Il�,H���Sc�ǷrTX���3�p{��2j���|�?�_���l^F�Zsv�͜�^�e m��xE7rob�%;�z�:4����� >���d��}(����Cs������a�Dⴖ��Z�>��N1�TX{��_�5OȾ�4�ں -�;Fn�� E�l�3��A����1:�G�����ö%'᤟8|��H����	M�"����"�����[�W�|�U�����:<��7i�� ������h.B���6oaV���R������{dXwv�r�5fg7�	�����ʈ#�B��'<��}��fJ%)��Wy���/iF}�Xa�o$�?�K�v�h�t�{i8�O~�1����J�<rL=���Z��]h�a^Y�I�:c�'��I�5G��t��2�z�U�ӊS��D��拢W~E��7��m�Y���ATh��*�.T۸�����(6-w�D?�f6�GT����EwbXE���JwJs�"9#b��������m�����Y7)$��]�w-��0Z/�j*��׳�Zp�JXi�C(���k��؎�h��F�U���*!��ܑ?K��7���ߥD�~Jk�'Nb_,I$j��>�>��)f��� ��%��ܽ�	.������ �?r�Y�h�k��SkL�sc�Y:�x�pp���sG�)zI��6#-��:5Ʈ�:z��]c���%Z�%�M��N��1��F�U��������!u~���7�F��]nʊ]A�<GvHvD���di�ю���� �g���]SP4#����GrEqR֒����$m��@	���v��<o�j��d��ʱ���'l��������������fw�e(+���C�^��[!�f�<_����;!)��� 0|�E%*-au�6��In�������;w*���$�y��FJ�׌E^�e��j�@q�M�k����-(��y+����oP��c�pr�J������_/Yٗ��#��R��G0�`���H�M�	ݪ���,0Sg'���o�����U΢DRvu {�Q�x�r��*�EA��[ik�1�����O����S�On<wo�u'��eN�
�e�MKd
���UAT��X�D�'��4a{�s��:"v�1@�EJ��nkT;�ez� ^lR�uW����>Ȫs�`o��s�E��\�"�M�p�]e�xoy�ƥ��߹���?��OQY� )��oM�;��>��I������U�c����{�	h��OV�� Ħj���N�÷����BR�(�;�1�������ψ�e�H�����������b����s�_�i�}}H�C�/�)!Uo�y"��X��"JA��"��?Ԅ���%�V,�Dڲ�~ �'@�Ƣ��Ԛ���M�7F���b�Q��Z��	�G�j>L�fd�8�g�w�ȡ+�������Ƨ�Q��s*�,z�@=����c�K Ϝk�9���K�_�כW��ӛ<��������s��lle��t�ٝA.Y��Vi����0ٛ�`e��O��q	����mrG�i�M"+�,d��_9=r?Ky,߅��G`y�%��*<{�11�[{E�uMK��U�RM(�˅^EF�W�)��0�rWӷ%m��ޅP�3$���_�����!䕄�-A���aFUd�����B��h�p�y���,#��n5J7X.�-�hb��B@�6u�/�ƮY8yr�P�aD32�2S�� W����(��R�#����Q��0�2�?"�@�&G�HB��<O�t�:B;Fv��^y/f(�6&�
�v��[64�f(	�%!����O��Yƣ#�2q}����8Th��(ͱ��d1�X~Bu�'~���,��9���}8_��V�4�k$�o���R�����&���e��,V�E�7��I�Xl�*��J���/�}�m�U�|Xe@d�0�ڍSO�
�׃:a4ҷ�}qζ꾃�5��x���#sW�"r��z�Ɣ ch6��=�b@�Qc��M��a>��[sQrɭEF��|��"@o���
�!�P��b�W��a��ҡxaU�h��n��G6�3Yp��ӷ��{�x~�`�LE�y�A�D�\*��?�v�\������*ƚP{H��Sc��(!w�R��6�S�;�2RSיE����+�n��<�L ��T�]N�7E؊�|!���;c�Wu�{xO���^#z�_Kw�^��&7Ckj���3|^J��e&��]5Q������9�lE�v?�+_zD�j�,nS���n��T��7@W����{.<���4�40�s+K�k0?+HY��Cœ!7x��+-Ѱ�X1�=�{v1��Q�~�%>����zrw<6��+��� 6���]ܟϫ�y�D�JZ��8ZLz�Nۭ�^@��ڠ��/��C�/�t���qD,w5ۯ���Qh���ɗ��~�߼[m�*�nzd� ���J-�` QX<5ou�W��e���6_�D.�_���?!/�0~*2�!�h�~���6�ʱ��4F�N[`����O��s)���q��P���Lfr���<.E�v8Y��z,� drdo�K���*�}�Z���4c1��qM.���@ۏ��M�\9�)c�f(|r+��_ �1�+�X�¤����U�h7pvxH+�	���?��	�|���p��H�(2���=�6�]e��e.C�'����B�Q(�~�;�oâH��v8�缠�l��Jmx9i*��9�2_�H�F?��2��W1Q�L�
��FRO� ���.s�p� �K���x�:�-vp���ޕr�HH��YJL�'��Q+R���
)&��t�3}ހ����]U/�CE�T�l@�'+����ttº��)l�+�1n�}n��W6>1 s.:� ����+�s�V9����i���B�N��vr�X-��%�n�c8�^&��tO�ZIJw�/]z0��1��X?SZD�c�ĸZ$�R�!7�
ǯ��N�X��r��~7�|+�JgyI�L}��ͪ:z�A-���g��V`IT4�V	';�XW�=��I�NhD�Cg+���/��x�'ھ�;ٓ��6i:���"g���9AX��T�������B�,���һ���p���	z�I�z��a���7���JwA��]L��;�_4�VP�R�2m&�=%"��t��@�Y�'��Y�Y���2�Bah.�i��ޥhTi_�'�� ��Ӳv��nE��:��חLE���I�4�sM��~D�ڊ#��p����ֈ�i�!ؗ�T��j]z,1O~G�׫Pn�5t����mm�"˜�r��^�W�̓��/w�����[���5��}��������䭺İ����㋿c���.��WQ��U~����1ZXfч�����?��� �f�j�F�]ICm�����^�K,"�W���p�=��G��n�[��-�������	�.��:L9Po �-�h&`zQ!��⌺��a@ο�6����<U�
��#��CR���}���ŠnM�im8���9�H��Y���2s^��b�G�.����wfZ6o4c1>�\*_�Q?��P��� V,�Z�K�����z.p8���D<-�S�4�e�!'�f]�b"13>�����<W���Z��;�����g�-��e�P���vA�ҒѲX��b0x�'&�m�@_f;�,e��B_m�l��5�����1۠�4�pmGS�
�M�q���a��33NDY��K6}���U��$���j��	�S"ъL�f��~48]�6����OZ��}HЭ�5�U���H-���zֈ^�@��ِ�~KɘeaNN-��w����2bi��a�"$"�t��8
���-xFpF}:g�~ŷ�[�b�0L�Jm���L�^�B��ܙ���C���1�1��-�$S�+�"�a�Y|k��Gc=�A�/�u_���k\��.�;蔰�C�h���z��sv���a�h0.Up{�ne�BY7�B�Qd(ng Ş���R�<�O��Љ�ŅD)u�U�Ĵ�ꎀ�_�������ViDۛ��+�2��#O ��5����`����&�n��kꝔ�_M�գ�!X��OTj䔣���#���o�2 P�ʰ,�|&�	��q�>�]�C�8d�'��>A����.6�b8�Z��N�b�j�}�<�X;_��8�`������	bs[794״im�΄|�Q�m}�Pa���ۆ���������y�ݷ�V�� ,T�z�5U�bx�k3j;��knl�J�5���`;�#w��Hk���M�S���\�߰��O�n����?{�y����o�a�ұj�L:`�	���T��z�J~�(>էf�5غ�?�SΚ��A����u�9�!s=��Q�����,���d�b��JP��e7�kΕ�s���w��J��{-�~��Ә���˯�lb܉c�O
8��5V��}a���7}�B���I���2��:�f
|�%�.;.H}�8O�B�ZPw�IR�2�p ��w�ov��L{�}w6�&s͖)RU���Su�P���z�-��iC�������ܒo4N�R7e��S�rSd�x����5�jn9Vk���6��P�A��rQ����	�O%���%�=w����˕�סR��㡸��;F����,h���?���'^#�fY��H)~�îm���r9��^�l�a
�:���O�U���C�8�&�Ј�B��=������)!7Wi��J�m�Von�2
�� ���l�^���M�-���a�Q���Y8$UG$�u�y��\��<EZ�+FI1hߌZ�n8�=]����,�y� ����}�ۡ1���?��`��~��ПZ������������q�D��;����k���̄5��G�k��<�k�l���@���MFdh�pt���� ٓ�z����M"�.���.e��[>@�a�)FMm�q�/(�A)��f���\T���ge�a�z#��LD�Nt$_8,=i;� �w~�`^G~���1��,���ĺ� �˯f� ��*po'	�YN���~>�A���:�Y?���^>f��kQ��/5�����c[��p��vM��V�$�'>�5<�����%���5� x6hU�e�r5@B,��Iҳ�M[�bCa�Aw�xMn?=Toxf,A(���끀��#_��H��G��� [թ�p��8����X}��fW^�S.�d�ȶj=��4����r����n��m=��kVnL�݇)������R}����b�	��.U0ϙ�ݤb��wϼ&�h��e��I��B��uZ��u��o�䇃��^�B�Iz��\�+�rVnW=K�7��R�@�	<�|M(��3˽8��&�Y�(���<�H��0߇���S�	��d�LF����w�ίϦŷ/�a����vD���Jj*�~���K��1����2Ԃ��􀃘�h�(����TJzs��%�;]M=����?�c��ʑl���_�A+��� ~tI!�|$c�?%�!��Ɍ�>`5�7�����RD�_�u�I}ט��5�T�R��ܑ��ya,���w:�a0T�b�g���$f�v�6Q^�/�����ɽ'I�S�D>��0ːNUl��{�3�EZ�|ֺi]��0�$�dUA���������16�����Ҡ=J�M���5�.�V���1�/��H6���������Қ��@zffro4V$s��~�0o�bh�GL�K+�>�}j	$JϰPuȋ��z'<�z����R��ՠ�c�=��#��N󠙷 J�ȑM��F
L�y���%g1p
H擌v��F�5pQ-+0��>���("�sy�?�j��W蕏��C��p���i�%�P��E��f�C��s����T�@���4O�_stf��׾������|d������q���#���ĝ8W�6y�^�q����m�ӡڴ�J���Wy2�+uo�C?�؁�"Z��ZyxI�t����}�}R5�� �e��x��v&�>�����}󣹷��}
�x�I�'м��LO��C�pB����5;��]�&E��'�t0nөɶ���-��\��T���х2gR��V)�J)n:�:�W�?T��42���`�;���%v�$8�"��k"�o��b����G���	dV?�;W�R >�e�A&������>���ݿ֨M�>Ub٢q�!���4e��q/�|}�,�Ir��ܘ6&º���c`w�\ENu�Ĵ?��^D���Gcj�)��FHs���y�����^�v�����Ke,˗5��}K���}7���`�Fs��
��$V/k}B,O��R�$�<	.G!�?�������+#\K��O�r���i�5�M a