XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A��W��iw����~fn7'���뙑�B���3��U&�i䨩�I����>kF�E�7I�?D��k��+������?���Q���1���#�_drg常X�����2�5#XZ�q�VxȀ�s£�Ae@2	��]n��L['�ά����3����Gj�o�#ۉ�8.z��W�[�S؃Q�b�%�UOGe�B���?
����l����� ���̀4�Ax�j�#�L�;pAzV,s���&���k��I���]<�pAr�8���]�νd�Ӌ$�;w��-�+�����ugȍ�B.�0�|N��R���>ڥ�gx��8���΀�f�_H�o�Iy�٩\48��f~ޣʂ���پ�$�Z�t�~�_(�~�础e�$]x� J�*E4��S�����1��|�f5�'E'��G}d�.AV=Rݣ;n�ӎ�^}%��" � �[�80�Q�ik��x(�������M�t�Gf�:ԩa��	79��C�#��p��*���\ˢ�_9�-D�߮�-���+~�Ie�]"��G�ĕ`G�B��c"11�v@��}7E�\k&�Ճj��D(5iFof4����#� �r�]0�� �`�B1�T~�.�B�G��t��`�g*A$�\�����\�s�n��
	DZH�&9� |m��3X#���q��S��1�?ZQ��*Y��״hO��L7x���?���\9%�N�(���"%̥��ݰ:�O� b�PJG;BV�a,ꩫ�h֨��:Y?ʌ�XlxVHYEB    1b65     a80T��R�CEum���r�1�Š|Gyޒ����޹SS!��*@BC-\�9=���L$�Ԋ��f�mnE|��2�̇��&e��[o�9�c	|��U�sւw���V�-eأUg��Y���c3װZ�������/fM[�=��0��ugo��Մ֥�`�VA�H1�T��dsjm�F�I������]���_��<Μ�]{Q��^�C��H:�R���iʷdm��gӻ8w���/���'�ʵ�Ai�+`X
���]���Ca*���)!p���;5P���ߺ�B�g ����"���C��tPn���ؽ#��p�a�z#}(6�~��1I��H�S��U���2��R��`ҭ��@v�������o�g���ݹ)�	�-Rw0�>�����dXeu��[)�ᢖ]��B1C3�%��d
1�6+�����g�9��.tڡ�j�� p��j�iB������vK��M:��Pf���f4�{b��sܦ�����4��K��`�vW'X�*?�_��wS��%/X7�(��9(@�-�ۑ�ʶx������E(���.��K�~�2�
�M��F쟽R6T�/ĜQ!�ɮ���yxZq*����$%\a�՛D�#Э":,֖�r�u��,�s����>Z��}~zҥ�g�B6�z-F�P���͂IZX<8c���gr��i�m�O�$�Ȼ;p���#c�9��\���N���*'��
X��?$4�pb�b=��b�i3������ZS�	�s�>�޺y7�\-h|����k�����ib*/�"5v��Y{�&(�I�B����y�2=�N���{6�r\��m�_;,���J��J22.�y�vV"Om(�;z��:�������J
�Jlq���^�p�}r" <�,���n�p&���"Ǥ�  �$����I�=�lX0"|�{���
���^�pS����|�)�+#"q��!������(,و<�^n�?�b��q߼A��9�Pu��h�`u�)Ft�����mk0�k<È\!�V�e�ƶ w+��G�����	>�� t��y\������rїM-�����}�EX�O�kw�n��G4A��hli�9��ϛKDhah{��0����q!]EWoi�%��E��;w�)S�X��{�U'��������oW92)�Y(6�����㸓h�p�+m�Z���G��At����&Q��a�K5��S�7<�W�=�$��Vx���]	 o��FX˘އ㘳�����l'��@�o��b���9H���Q}+(EE�l\s�TN۳�ڭ���LzeI�H9�@՟�cwBʊ�B�{��W��?��(A��A�X(�6�I�J��$ W���E���t�m!�Ա�'`w�k�w��j����8�~��fn=�'�&�|��Yl�	���O��*+�]U���	��y����$�n6^��P1ƇQ�D�Bd���G�_}uC;/����PO���A���T�I-�K�w�s�D��
���e#���Ye&ҁBD�r)dm$<4�;�_f�e�i�c��zZC�kZ>��N�Q��2��j��X�J�_�w�[x#ל����i���{���F��8�@,Jf#G�+zn^�)�sB��07���w���X&����5	$<����A�.g�ë�E��p�DM�U���,b�T%���n�S�ڔ����.�,�@~�.���(F˸�BGy=ŉ_GM�ZFIU�;����`a^<꺫�Ŷ���U�̊�-��/��=�@�`L���#5@�1�lX�3����謽.�X��Vw�8ht�DP{OU�]���c��0�ْ4U	��腅����QXt�>~�Ĕ	rF+b�x���+_���@O�-I@�d����`��5��d�}d)��Hq�:�5i��T�>LrY�4B:��u���P�!5�D��n��Lr��1�'��2ua�?n�j�W}�l=�$��qM*��m��p�h���YB��$�\I+�o�o��<���2��sNnc��0U�M�e�E���^BF��7E�yJ�c����\J'�Ӿ��K1wJ�ʿ�����ye�)��V�-�L86��L=<�n����W�xHS�K#�w4c7���*����g@b��4���/�40,���,�c͓�����<hP�:��p���{x
d�4ɨ5o6�����
;*|I符I��[��6ߋ�S5�C恔�OG����P/�X&�ߍ�k��t�3�!Ao򿨟?cٗ��U����O�����ꭢy����-�v3u��a��V��k��M�:�cK���8�}3]*��u"�����X+�M]s}���8I��&; ��s�^4�&�{�Ԛ2��#:a]9��6|�fA�����{��>�ե�dV�F�l���t���wؔ�U�C��~����	�9�~b�]v�	ŷ�����k�J�z�B�Z��oOl���l7�
��+�k�*~߈\�ɜi���p�u,��4���nk��-�r,q?��)T$�A"��!��0~EL9ӛ�X@���l3r<�pRJ�"��VNɘ�I�x��N��K�٣��ϐӍ<L�RD�Qx@���n��%C�P�#���<��&������ �SR'�8{�0�9�N�
T�����b���/�6��e).��M~Z�J���ퟸu��ctv1'�3�ú��0�'�����'7j�f�E���FH��v�W��`0�2KL��