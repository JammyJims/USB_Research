XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��md�.�h���H�q;J�d�짴!3H�
l�S�*Fx	aH��A�Ɂ�A����0J���n���_�mGl�x��h?��}�kv��0g%�	�Ї�-ߝu�Mɍ���b��7�dH�J{�͇3(u�?k�4��kE��� �{I����Z��d��A�`��5(�+]��K��;k�+�+[��b��j7�|H�y�W�sل̛�q*R=���bFX�-���܂==�����U����P"��#������yP�1�^��1��� 1�g�an`̖S�	�цXR:ʐ��u�����z��EY壈��+r�T�w�'�Xo�yV��x?¿ꭨt�s����媰nd��y��,�ƌ۲�!������z�T�y�t+� 7��2��"���T�X�1j9�y��s��R�\]���.��0R���~r��h)
"l�B��꺥
*�mǍ�e�ʷ1��r&��wf�i*��-$����,Wi��k-_�x�QV�����I�v��+�l�Tؙ�c57�q�
t������V?-#�mc��e��Q�6�|g)�ۉ-z�xV��,N���H�ѱ�d�g���	d��'����vG�X�q�X�&
҃1o�7���%����q�A}Lj���[����I^`:?fP�g�'�8z�(E=G"��������@,ڙl**'h;��r�sRk��!9�N/�u({۠�����Њdg�4�>���(�L���&�����R�Q�2��f�ٳv�d-�&?mF�ı��t�-���&9XlxVHYEB    9bf8    1d10E�8��k*sP�|z�0��L�x�� �ϖ+� SC�O��������BK�m]���R��Ub�#7s�o�|��N�m�%�ҧ6�zc+ߵ��������nZ�["��d:����1���1�޹b����Sv0�s�'�Ex&��1�k�퓉��]
�F�3���QY��\@H�iR6�i�U�x���q��13�"��Y�(q9Ű���W����*�R��!P�Qy! t�l) ��0ɘ:�C�*�^}��q1EN^ >����p�-0�3F�)��	[�t3Xf-��U�A,�����(�EV���B��=·0ʨ�Ѐ*^��p��ؕ~q%��d|�?/yW�0M�K�����m-���\���r#:�G�Ec�}�J��Vw��S�~V�oaJǴ����v2����00D[
g�t{�>��j��}Oʄ6�tA8C��AnL��-Ȏ�@{���9�nK�`ljPb�瀬�~��)$�Z���g�@���>5�e���w�v0�L�b-�U�k�ֻX�b��CU}�=���@�BF�B�})�c(=G�^7������)�����c�� ���.3�3�2n5�f���]��IU1�F��p��k³d�`!c�Q�]��e�*��]�����p��j�y��ݼ��nw������UH�GnQ����{c-�?n �B��eʄ:��~d��I���gG�J]Y��"�4r��;E�X/�}����z�7�L�b�R	�BD��Boz3$��9#�;�W��	~$&(#��(�	hQ�bL\�-�ƾ���N�?1�v龱���mJN>�~�ZN�@AO6#L�4_����l�o]��O�,087����i�����;y����Uq�Ɵ�O��D~�2监�F=ڎ&S
W[��#�`��F>"��a�ٙ����K^��ћ&d:f�bwx��l��쒣hN(0l��t�C;|��=����Tb��O���/�'Y�E��C���ڜ�9�
^oBaV0Y���o��"k��4�f�nx��@^Q�	 �^���"���1�[Q�@�����Ww`��,��DK΢��I�X9�	�_��WX#Zn��]��b�T�)���}�U��v��[��IA�����Q���Cj�{�8b����1��d=$��,�Q���jPP��Og�@�|�ނH����k��:�6*k����,�jh����oI����h�H��苕����9G�ߏķ
4ᯄǿZ�^�4{��=��G��N��������B��P�(�`�@����0Wr�V���L��`�� ��3S��	.-��F�!a�K
\7������j1w�m� b�`˥5/��9)xR���Z�Bi	�����7��݂����"H4R�ƹJ�'x�����fv��Z�t)��~�yE���I�"s�O6�h��F�E�A�����"��>ju$f7����P�`'K^P]��P����N�Hr������G�ǡ�_/C����zرX"g����#�8�_��f��}\�z��P����'x�^'7O�"UĈ���]u$˚�C����f��Z�4��fM
�����KZ�P�r��o�:�K��]�Y����<���E����41O�-�nr��z�����]���������B� HM�Y��i�i�@U�ק}��R���v��*�j�D[�;�oM�*.��k�:P\��=V���[s��������ު!��u�P�/l(f�[3N+>��ڞ	)��X铦��n
W�:�	Ux�$+�6�d��im:>�t�$y_$ڀ˼[A�L�i�^��� �t]���Kԥ�� wE8�f����5�˫X��x[ڜ�k���]���L�P�����X������e:��V3Ax!�ʊ@�I���5�;��:"�9�V�a���]e����a�^���������}�t��T����M���rjЇ��u&��f5�/p�BŸS�O���LOi5ÚEK^r�O�����P+>-�{d�2���/��?:eI�2}�Ⱥ���:����wimz�0�Ǖe�8����x� 0�5�J����~9��I�Ig�$7 ������RF{Zr.]�8Y%��Q,%�:
c[�XQ�\�vVrh@���e�,(JS������O���S� �!�ԑy8�ڢ+�B9pc�c��>�W��/�t�)4<�^���H��`��#�W����2�����܎�n���v�u�/[�q���BqW��Y@��7mo�|:fH�ߐI�[VP؝���r=��a l��6��Ӌ�P���~t�ކ�dNQ;�.3C�F��7ye1�cƕт�|@�����c�inV�Ȳq��awL�M|q^��L}���-i�������"�0�'���kj���B���Jٞ��'���;i�r5��p��0R��1��(?���zU�w���Դ���'�3�zJ<R�x>����Tx�����6cn�H��;��V1M�p���ѣc��0_����DV��)a�5똘Ҋ�`bis��L�)vo��#,x98+mdm=��1Ѝ��p3?����P� %3F�b��
������]��@� E�qq��P��V����da5�
c��s����E�ד%��\n|K���,v�';I*TĽ��`����ҨS�^|��Ě�KN"�YJ�ܶ`�UΏ�� ��*��5�Ath�c�P�4��!)�$�b���-��kNS ��Co|�QD4��6:R�±QQ���㉈�c��c��2��|��8�s����o�vE��W��6��,��0���\�H:�z�h�N0��+ ��~Ø,;��􄄮*H7Ҝ.��C��v�؅����.,�=����Xi쁚9�h�Z#_ʗQ�l�~��ܽ���� 3l�q��� \���� &��K��TE�<���=�q���<���Wg�
��~��X� �9�6}Nּ7u�����p�cw�	.��F5�#X�9���x{z21��[����QS�l,tq-3��"b���@��ۈ�) T�G.��R���-���`�f�!�����+��t�����G����Y�lВ�O�pOj���Ey-�]��g��y�D�hv�������r�Np
��6+[�Vi�31F�rKx�I�5�.wBZ��>�Q��HN:�qO�>k����"wCUX��{�՚���_j�W����)`��w�#�G�E����ҵ���n�p!�y��0��޽<n��E����h�5�>o-A������`�˜?�&RY��D�s�� �pˊ�l�Ze.l��GP�K/#,�Ow@/#�m����-�U��ogD)������\�aR�� V����ۉro+���GjE�-��`�;G�xX��������;$^�dā;N��&uWqM�X�v��f.L��[��g�Z���n�.7���f^T��d�au��}��%���2�%��n��<��@�v����J�����2k�WZ�vErD=6�5��w��@4Ř��5��򽄒�j�п]Cѕ��B$.� ��������5aǝT��@Jդ����A7IR��L������6,��� �3:�-y�N<OU���E�������7T�z�L��B�V[3�@[�Jtl�4k�BPlo��M�v���-ݵ2��@��%n�! �9<��2_14������t���]f����%��$�|B��1�J,� D\L�,�!1���Ix�I'On��eL���Ҿ��ސ����!�<��\ڨ��2��5YI<e��:�˵b�PH��v"�Or;H�|�~�*��l�67&�J����p�H��!��4�zh%P܎`�c`�>e������nU\�ŊAM!&Iy���;�x��Ϊ��>��:7Dw�UD4��.�49�hRC��Ƈ��X�׸��F��nie�y��Y[ϩ�����2��������i�	)R���W��924c�||���[�����?�9.^���3�0�h�a���,�?������)%���6�C՞�W1�M%}\��kW3�t&5/-����� @����f� ���9;�0��z�F�~�	3�j`�o�PD��Ƭm����=>�类-ҕ�L�/:�A�1QD1�T���<2�%����!4������վgs�����SU��m�yJ{,�䈶�L��M?b��@�W?p� ��5�)�&�wN�t��5��0�K�W͵�!��#W��uQ&�S���;�-'�ض�;�L�W\	7^��Z��x�}�ߊ�F��."�7��#�W�ٌ�Lu 4�w���\}֝}x�oY�$�:��싓#U-��2�36S���Oƅ�W��7�=Gv�Ʌ~f,o�q�Mķ` ��(q�+�4��u�6���ǝ���*\Η'{4Rٚ�8�	eqNy�׵�B���W�&+���o1:|V�]�?�x���<j���>y\�X�0_~�n��w�(+�8�-�$]}m�q={"��������U���3���Ϧ��]۪'��$]��������==hg��W6�B��'��ۯX�N{Cm12�?�����A���������KY	TWeD%o�J����2*3`\� �q
�Ga|{^4�YjB��U;Y�rF��sTn��0�M�\�T� T���$�hH�W-�_Qrӥ�5��I!)�R�M=5m�����GV6ܻe�˯mFX���h��;��5EsUUW�P�^����W��IK�g���1r�F��*�?��}������@QIf_��@SY\A#�V`Z�1�P�����yIl�#h�of3���/�j�&�"K�:�8��L��p-Z��w,�4?ᖺ��]��C�͂�0)\�������zo���}"�˽���sp��j'�7���Pw��Y��l%�'�O����1?���c��a8یK��ք���3�r'hԙ@"����C;Vݶy`x�el�V��R�?�0z��Ͳ�ְ����R!��R1Q���W=�Ot���l
�[Go�](A4g�3D��'�-�SI�VM3Į^�A��( n�[��-��҇��K��ο���.����
`/�DlѢC��9D���r�ӱl��d��mL���V'��B�����救۔J�|�)���9�����5�"�4�'b���+��
��l����fJa�!a�.v/���0��+L���K?��`�=�⧌���ھ6}(�~�D�0��09$�,w:ҷ6�3ǔ�5�ŧ%s�u�Co���Bc�ci�	
k�:��Dp��*�ЃtL��}��2wt�If�a��)ޚI�>�J��D��R!�3���
��
8�R�	�>㡽תѓ���+�痦�����ˀ����=N�+�A7���N��D�p�?�^s1B ~��_}~3�b����ŷ�v�G�9�s�`�dN��K~�+�,L�!G���.C��}Û&�q���`�=U����釯*S�1��
�� ���!M�����؜<�,���O���X�R���� ~ �Umo�p!�d��ᮦ�@��H&�ON�f�����`֍v���2L$�=�}��VF_��N�x���	�L�!�)��&:��G����˧׽2���0A@�Vl�w�6}�3����%��˅`�It��^�Fc�'�r73���u���GAk���	f���n	���NgZ_�A�k�?l��(�<4Jj���x�0�r�a�V�޹����a�� ��ј��/����u\tX�X`Z���3���>��.��*��NN������Ac�1C8wG6���7�ѐ&�i��H�� ,���2�dL5��`��Г�S=�OK�ɍ���n������o�4���p�ڛHQ�&�U��}��9ݛ8�y���F�:�൱C%�k/?��,6<J4}�D(�l���׎�a�!A�_�Qʸ=���
_���>��(��ګ'���W�-,�}�泺�f"l���'��v�I�n���.�ֺv�ب��(�OA�+���gt˹�a9,h(�� �C8p�@���������>2��KI���b o����y$���<��n�WZbN"�^{��R�R͛q:��P4 bV":R�fkD�'"�yP4���M�|S��иs\-���������1�뺣E�	6U���.ei{L����,��OX��[U,^vj��`���#V��������,h	?��tL��M�B�#C��^b���g><<
;����eH_��߇��
ꋘ��mPjD<��s����A�@Y��M��L�+I���Α#��ធ�5��(����'	y����&�d�ן��f�N�d1'����%�������u�_�r�<��v�L��"�9B�Bz��{� �N��Veƃ_9��$��	�FqڀU��ݰdiIܱ��_粃aa9�p2Ἐ�1I4���\�xo�p�^|�dl%��<t��p�;].I��}�q�`�}�z���ĥ��]'Q"��&8f=�����~1*��&��~p���+��L~'����a�c���SH�/㖐�ّ�4t6����Ҭ��G�����n6"޽�=��l/�s���u��a����w���؄�T����ݓ�6��`�m����[��
��W<�
׮�ΝV�V0�Q슔M%X���� ���:^�o�<�J��g�"�����+�0�}
�σ���G�@�]�>B=v���t�^���F4qN�l�.� ����4�@P��/i�Z�p�vu�EBG����E���;Qq�]3t8�"aX�l�
T'�`-�Z�S�y6g4�65�u`�F:u���sE�i�KL4��Ga� ����~��
�o���"j:�VF� 5-��q��:���~m��m���O-�.�z*�+�Ƶn<�1u �X�g�߬^�\QiuC��E>A�����&VN��	̹��}o�a�5nK���Ƚ7N
���H���sضv���x)�	��:r��#�v�D(�~F���l� �1M���#wY6��3G�s*n���^cAVfEnк��Ò��� ���FpO��Lh�F�T���(	�^;
�S��;u�)y5c���L$*ʭ��mo<�$�?:�Np{��M�~�% �����WWQ��PN�|����-\��Är=� h^@�,X�v�L*5�rc�q^vE�HG�?D~��� ��M^�be pї��r���^&B\A47c�����ퟷ� C�R�1�ч/���X��?j���-�j6<�ߕ d��Yʦ@��T��-}S�/�q���F�e��d��=��a0v*�R0�6�� �}�����1�YE�������t��؊,��G+D��d �	8�� 4u�S��5��������V��������ei<�T�>N�9'9�{�8&|/˴