XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���'��7ѐί)i�8�~�#�P�=Q-�ǳ`W��+o�� �		轐1)�<�DG��!�d<��/���`�$'��}E��%�m��j�y�6�.�+0,����fyc���	 ��^��+e[�����(޲�W�cs5���7�k���3n,��ܒf��``�`������0�*��O��6�B�PSo��1��q?��N`����� ^��/2Q'�nҊ,mTH�������Ew����� pf�U��U'��U=��nm%���,&�8?���i���}�}ǘ��U�f�0�r�< ��Ck�Z>����s�G?�Z��Nÿ8���|=c���mX �v ����XKHh�Wk^l�!�|��flT/H�|+gA���*.��+Ǫ8[I���$1-w��B�� ��6��
ۖ��or;��7F�tl[�}%�8��:--Z�=߼�0,5�UlGD�u��=-���!��>�(a9)@b���f�E�����o���c��-,���b=I"�!P�X���C��8���:�.)͉J��Hw�&�`��e�1�i�MƏ��V��%��#$(�d�:��> ۇ��c��K��~<��|���~��,i���܏�Q	�	��^�/���)��R�|���=D��MT1|���l��%�Z�ZN���*�aP.�H}��V�=�(�(~I���bB"��%+n��D�]o�;o�U�`�S�u�q(��0���=,��b_~�D/�A�ɕ�l}0XlxVHYEB    37cc     ca0p������k�)��B�py���@킲)�p_P����S��2���B���r籦םY�)�`��t4�ǭF�R�I�g�<W_��7�\��z�M�͆�h���P\�B�ӆ�]�FI���TM;�h�[�� r����Gh���_��� ��E軰֘V��Q�"�o<��2T�ܫ�+(w혻�^}�5+�-��J��G���K��"e���O�o_I��/2�T���b�
��C8��� *��-�a�aD�y��F�_%Y���Ö��=%�Ӡ�#�⊙�1�)E����"�c֖�ȼ6h��}����k�y�4�;wӑ<Gf^d�5(��=��Y�k���QW�P~�|`J��O��6�z��Pϛ�/�q����uH��+<�ߔ�`8嫫D>��`��(�Y�6 �ڂZl#u��v��ۛ�+�ňr��aoQ��zQ)�@ �dR0��L0ՌU\�L��<DD^q���Rr�r����]��o�b�˄.8q�m��	˽P�K��c{���0�q�Ї��$��4�s-RX9��޸�bW�AY� !d��"p����ߋ�w@��)�����(�*v'��F��l}�k|���i�$L�HOc����Sn�.�N��Ֆ�d^R֏�~���M0O����jE<K��.�:M���Q����ޭoMpJR���,�Z����Ɯ@�S��7On[@
��_�8Z�;�ǚ؅6� :�����k	�&�] �>��Xڏf�Z�ń,8[��q'>��(j#����"��Vڭ�K(]<u�թDyCv�$����h���v�΋��럙�*!�����i�hr
>�=r�kp�Y��I�n��A9�Z�n����	Oa�3#�G� U6��i��=�lW�=h4ĵ?�aR������K�����Y���/ ����Ր�� �
�ܿk��ӷ�;6��)�V��cl9t���hBRWϙ)�')��aC�X�nG�)L�G+I�Pe9ͻ���!Cɜ��~t��puf��z{����iŤ��ٹ�nN`\�|g��J��?�����ѹ�J{~��6��d2�G��j췜�4M�wϘ�KB*�;	&�Ǹ�{uI���n�b�����o
��e0p��I	�aՊL`,�ELA�� ��ޯ��<y�/7r��LW"�D>CˏY�8�m_0PY�d!'���_'Uг$<>=�"dX����3��J���T�����nQGFn0�H-s�n��*i�_�ˡlf�j&�r�Y�|A��\Aq�,䝤�>+��J�
E}u�W�:S]�}�4����>��y�%�69�5�@�5"�xd���_z,�`�l��^u���w��*�[s�(��V�g0��@z� @\e��:���Z��Z�ES-��xP�&3o˨�8ט ��^@�J����+�x�Bt�O�����q�̂������̣<��ONh`���ؿܼ�6�����
V��������gU�T]��%���~������EH{���^���#c �"q�ztJr�^��O�������sՈ4��l�Q	�6�!��΋=�(v��	c��Ԋ̱�0���`O���İ 8ʣHt� �� ׽:���W�yBuz�Jf�Q�n�����
/_:����/��o��T��2�@'�v��L=8���<��"VE7�؇������J�'�%��� ��������ƨf��<'�F�=�Z(z�k�{�o
jA����L��t���	V�Ҟ��������J�b"�fy��J�L-���,ꐊ ��H�9�l0���'ȗ.�V���W �&��s�N�d~���f���g�ݖ�*y��R�ڦU]\���T�*��ٿgT��+=A���Z����"�����x򙀆�.��ͩ<�i�_QerWr�L//򌓡������FMК�Y�\}4���%��L�$��ٱ�z�X�Փ�o?^����j<�bX��U=_)�6$�h�&-k�����[�s��Y��
J��&�3.z�X��b�\[��ٟ!]�.�3��ܪ�d�kss�����#��ۛE�O��FSS�%�"�:�ջ�J�@��O������k�?�ƚ`t�GT;�P����ƒh���`�eMas�1�)���~�xia=MP�,��]��J׌^mNW,�n��dF�p��P^$��ᑇ~a�V��"`A=�N�p��z�Y�RE<]n���K.&rFhw"�.Cɩ��=?��YBF����my�����r�貄�}�K,�M�=ē��2J�m�Ks+�qu�r��q;�wY�4$�&B l���$yg���xpH� :Hi��_�ֿE��5|h�S}!Mk�n�X5�Ϫl1����9εչr�0n:m=�dV685O�,�`~���ZR����x�.[9���w��fx�J��a@T/	Z���sc��#������.�r�Jc������)��:��0h7�ܦ�4�a܆�����y����Ř�C3}�Ab�C���SI[�ɋn'�Ӎ�g��K�Y�N����i%qd�3L�w�S�`dE+�C�-�I��R1a��9(��,w�J�ǆ.��|�,bc�r|�uq��%]�hW'�e���z"���L(�@K�L�H��R�܉�(�a2s��0��`�z_�6!D�:��?߅a��55c�oM��N�ۺ��z1i}�9�������zJ����B�y�D��d�D��&4zH�L|p�)��X��.�7���B��s(ja�� �6�5;s���JK���Į����#�4]��"OI�����	����(�7���}���J�LWAM��|7�2?�N{a�dDǟN�� t�ގ�'�M[�WB,��ub{����k���?ԺD����x�~k�쾐��K��hÑ<u3��Dt$? ����wB_�A�SLKA	Ws>�y��#����}���V��G�<�靣�7���V=�������}��yu]�^�|]L��6�B��I""O��N�#�I¶�RAb���sv�Rj����i�(��\�umQ�Nm�#XE֘f�fXNXLv�k[D)pK,��qRw�>��FK���:��j�=���垚�9u;����D܈E��C�%�)��y�H��"Qs7���m�Wv�Υ^Y���KJoN~$!K�93\4���6��+�,ުǻۧ�q%�