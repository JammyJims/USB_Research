XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&0�m1��ݷ ��%����77K���d�,�n�4��;��;�^h�d�|�h����ز���JJ)�T�z��r	��x!^nQK�	��������]/*��U�Qu�_h�9�8'�6*ֶޙR�Chx��w�:I#^�oxP��?���|�K˭�u�K�f԰P�y�����O(����&�2���$�u
[��K5���Lw$����]ǘӄ���ҧ>w��ZJ���}����%�����������J+���<c]�P����L	��I<IY�(�#:@1��cEt yG|����@	^qE��a�9�:!p"��	A�����jH���&�G2�]��|������L��Z6%�R\��_���YT�9�Y��u��b���F��Y1_�fg�"���(����m��w��������۾�qTa���m�S侀����7�$N�ߙB��-��rJ䴤yP4��A�����*�g�e��{������bT���,i��-(Z�Şx<�L���h�)	�GrV��u���C��.uvdy�o�+g�pYn�D<:"H������E,�zDm\��0���CUG[X^USW�<��8�G��I(Se/ !���FtZh�2�y��}3��'މmN�2�Mf������r�/���6S`l�nL<��k��-��Z�|u&��Ԇ��c�t<&Ý*Q���[� \��	�Á�W`�_m��ɩ	��]Y|�j���fm�ߨ�cQd�k6I۬�	�E��XlxVHYEB    2ffc     d00�H,�rq��ͼ ��k��8���=��Z��oc��.�%#�Sۊ����	��5�0楧1�aoצ�<6���� X�G.
�n=P5zrm��3x_�du*�XeM7�K��˳�7������ 8�!��	e��� �v>���kB��
��{|p���xƾ��2�: (�CCp�pw�ȡ ��h�HS6%��m�@�����⎪�mNw��ߎ9��'u�m �����N�����My�Mҿ��$��h��H�=,�a{y2:��KL�G�� 9�
��QF�`�N�V5�k�چ�=y`�� `��?*��E 3?�Fs����֍I��}5���dsyW �L��l_b��(K�ǂh�8c����%3~�o�΢�4��2�?!ޝ{��$�:yr�<>4;�AZ>)��B;�P�J�-#�ޘ�yy	-[Ɛ!0�8��͒�w43��A-�i$���ag��~)�2�'�C���� ���ɤs!=`F��k$X���a�w7ceg�;t�����I�ȸ��A���EP���K�b��Ӝ�ј�cBF�M#�б������<|*��D���s��V�;��4o��A*X�R6�#6������Y���@z�u����S�E�{;�GΡ�9қN����������u�zK5L݄<
�㚉i�RM�c�`�_��������jQx�(E��}n4؟]�D�u�1p�Z�#��N���:��9N6�i�����~q��xM��̮��>N�����R�J���~ ��1߂�󿵈��k<r��ٗ�y�!�
�;*�u���A���o0�:��4n_�����d��Q��d���v�A�Զ��k/2o	��[%��J���Z}g�f%�,�AI���n~�ܓ:zTnmXo�PnֽJu�o<�v'ǉ���A�VY�".ݮ���J.=]V���i�MT�*b׏4#~���L�>�7�u��g���fQ���!z/.��Vg�z0���3��G�{{�k&V�J&p�\��'޼�q���
��x/$�,�Z�-K^�|i��x�[g�Vf��L�59�ג��q���̳7DA��7��-3m�d) �B@����
�w�PC��,�� ���&���Q��͉ް�+&����@3qT�p��ߪ4,�Z�PK��j����포�n25&�3{�4�m����<�O@��tح|"%��y�:ޓ
��p�,�� ��Pb�)?1�JkLPLM��.
��*<�-�5�4����㹞}��sÈ:z�Qы�\��ܺ#SV`o�p�s��;��C-9nP�?F�c�}2{iSL}o���Z��}vӆ��ޢ�sM�~�ֺO�P�cc�����q��/6�nnS퀠/�l������h�#���J4(Z���V������,��p�'u}��L�^M��@8/���Qw?�dَu��q��:�t��J�ԅ�-|��w*�o�	G�z+���@~����+Zʞ�ʄS��	�qڟ��8,�|$*U�Ozmik��k��s�w�4愂�0���e� ePd+mXP���oA�dCB�������cj� ����}�z��[2�b��Q����+��9'@,��ld��s��V��Z������t	#_5ѻB�'�w�y[/�5���[��(��ȯ�<�6��^�\Y1ь���}�~x!-c�Va80D��5!Ĥ)?T�ن��3/�TX>Ӟ$��"lCArSP����������J�Hk��%Q�8�C�47R�]03���<��ز7�3
�PN����ieh4P�|LJ��w������@�E��5���G
tn�V��8.�_����Ư�N�7fDS��Ot�*��{9�f�!��婮�*b�:�P�T��/i�T�R-i� ���+a𝷕J�/M=n��{�k�*4�S7DDwyR=��' �ٖ�ۨ1��(���w@*�� ��p=`{S�e�ԕH��%��mU��]�����z�!�����Rp��.�<2}��e���TƁ��|�ُ3;�d:�R9\h
j�f�R��!�}�;�_� �Z����Ƌ<�|\Z���9 ����m)8Y&	����޳���35��i�	q7Hgdw��B��9OR�����n������P�1����*�H��|����ߢ�@�hyj~o4Q�swv�PB�����v����//e�*�� �0:��pg-����S��E���퐼U�.�����J�Z�[y�ɷUDi�m矛4�g��%P$O���&�^�����R��g��Ț۔��x�_gC��xҳ����&b6fq$��
�g�#&�����;��4dx�ys2��Y��'<��vs!�W�@>��D�H��^���/(�ُ���?1)aEC��Vr����E�Z�rNV]d-y{ey��k����`��@�	�;�:���Z9r�����׏~�W݃G�T��ڌ<fCZeG��dNl�'��| ����o�f�e�:�z�I�g�M�m|�i;��8���'~�21��	Rw��11#D�@��gQ��2l��s�Mp�k_��1���*^���F��u�4��C��O���䯱���G�a<���P���v?��F{����}r�MO�_V����U!��ZS�m1�V��!��Y S�AA@l�*����e�X�+��i,e�"|~�S��|�NYb(���M������m�7'\	�Q_��3�.%`U�k=�!L�2a{q9 ��a�Gӥ9��$&��N_+��'��y{J�V;�aIΠG��~�=��$قy�q�ۿL4���'2�_ar�m�	�������2���!���4�j�w^R�����"^��i���p
��w���}�Z��f��:]ّ������T���Bi��+�`�����J�}N?���ߎ�u�`�X�H$Q����'�~-�!�|�@�t]R 9w��@	9�,����GK��*#e����6Lo8w��bh�W^Y�o��L}�������l[�C���h&3�dly�FrUha�͎�⒌E�^P�e��ǫ�4�ڎ�,�ή�HPq��6������JR离Q;|����̊�<��d߀"�)~L�Mv���ryK���� W0�i<ub����/T:�(�D=H�� �������ՠ�^ f��|�6�D'm�o��N�I�X^,�>��.��]3v�������
f��<g���50�-=2�Bf��V�����������x`��j�)���Pt����/����&i�ߟo��J(+�%;O��^B�X��+�׳w�Ijnv��͢�����~-)Lh��`mcJ��bG�4�