XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u���{M��/J��|Ϛ?$�p+�
���%t���G1|�vZ�,
��v�%����U`M�[�y��� ymKg@Y�RX:����`U�x̣	�uJ����5��$(���im����[������!`�o]�8W{۽��_���P��'8%��߷�쨇*�O0�b���[��c���w�I��}/_��e�ʠ?u�6�TN6���2�r~�	��DW���5�i�H�}V�C�p��Qm�_-ˢa��9PS�Z�=A�]V��@�L?d\��hW����t�zyYJD(���T��g�m˪���ܿ��+G�iq�=�{܊ʲ&��4
?S�Z5_&�\	c����J�Y��5�=��S�z+��QX��i��r�nP�E��M�'�푱��ڂZ�XĀI��V��op� �s(l��i��&�	����h.	�Pі��?�ƹHѬ�#��g�������&��8������EAMZ��9��T*J+BHG�=\[�Ԋ"z?��Z�P_��wV�[7Pb�3g�`V�&.݀wH�Y4]#��R�̸)M%w�K�:��\�h��%��[
B��GY�a�+�*�E��b��ZpiA�h����.������]q�>杫8���%Н4�c��q�2Te�����TҼ����5;Ŧ}�rPt ���pKċR��'�7��}8�R�G^5`n�"�0��Ѝ��h�sz��z~�6���xL�S�?��!;��W��A8�+ic�^�����w�0�RL��%�'�\�"�XlxVHYEB    2c43     b80�š4:iֱ+9i���qT�lv�m�Ԏ�,���>r��C^FhђD�8NGM��
h�r���ݒ�n$wӉ�s>����1plU���p��s� ����)�<������C�T7+mVlfP��X0�Ĝ �9܎
;{l\����x�¾��_B��o���������U$����	\���t$�"�g@Y��I)��]<�R�x���iT�Պ�P3������XՓ�u��/�Ǖ�`�
��^�1��?���2}�V���ok��ɑEځ��X�F��`Q00�r8y�_ �⅜����Q��!�>��v_��bI�
��,!)�x�.P3 �Sm��1��d���un �t����+q�_�!�9�O�������\��R:�b���x˘\Z!��B�r�v�K�ɞt�Z��;�e�S� P\>�	�XH��#IS��+�(��Qڪ�����ݩ�_���7�c��0�b�F�
�,�XkHК��$��*0���B�o�)��s댩`��=��j��	7�ͯԖ��1�eT����{��E�@R�ol�0R��� ��tc�^�J&p�(���)mfZ�.p��h��$?�}S�e�]�#��p�<�V��vܒ�k]V���QAA]��`E������p�Qv�Ck��oD����ȫ�S�Q>���ˌX����i����|qYQ��B�eP�>�M"��B�M:��ϳ��}�A�[�YgNk<'$�o�λU4��V"�&5fk��S���j��Hb1[eLB�J���l�q����� ����s���8j��� �ab�ʲ��pܨ�n����E6�d�a1>>7��P�Jm74��>�>��%�"��l�ת��ʨfܒ��8eD��&]����{V}�n�M:�f?n3/�!��NռFD렼Atz�X��:{y ���js_��dkh����J
r�jF�-��.�9tl @A������'c5"��l�輵�o�I��;B>�t��T]r��a�;)�)[%5��z4����hu�%JG�	��S�UӇ�7c��2�.��S��e�ĥ�0��=�ƟV��K����yK���[?�L��2$����Q��y._$�,C��!<Oȸ���B(B+V��j�P�K��Ľ�q¾ �(ܷ  o��g���C��/+������-�,��/b;0�n�^I��	2ZW���Q���v<�I�l(١
:����()�'a����jH��U�e��g�L�8�����
z����`Ձ�����F�mԾԪF�|�lw�ڄ\�&$�D��
�����ٴPW�a�a����K�k�?���/w7����Q&��tfh�7���?S4hpJ��-��#��7A����h��i�u�y�,�q��'O�_��ҳ|�	�q�R	�74'2l��(X��kG`$�k�fn6����~Jr���4�V�~/����9g�W�X�v�Lp~8��#�-�M�c����_)�[.'���
�dKqT!��6��:��[F}T�,��vVMŨ']2�`���f0#j�b� �p�����%�����I_��^�4]J>'��U����wE �{P�� ��qN��s�����Z�r���2����o��xİ��G�!����'i$����̧J�ໍ��\ej�ɣԊazB����xV���al+pW��0����l���	"c2�B�[�^�{W�|�*F+85چ{+xT2~e0gW\պ$��ُ�żi���Ą�2Z7�l� }���I�d�� ��ur<^"%�t8���ܖ.�� `�s�&��t&�q���f��ؘl9�L���J��~��p\g���H��M�p����I��V|��(�O+�b�^�5��ze���[*���,&��KFz��=X9�����=�m�0���Ց)uQt9��g�@qo���j�:��(���E�{�`����EﲎDN�S��X7�$B���J]�N��0=�N��$!>[3/^�=;1�i���Пs�����0�@I,����;Dp
[�C�i	��B�#�;]1C���w#�:�_)�3��c�ˤ��o �~Y�̰��H[�֧]�����
���g�#-�Y5��n�qg����� L��"�s�
����c���%�=`������BW���$��=�x�3�SH�&��,�%�r��gGJ�8�	�`��z���z��������|�ʆծ��^�l��L�F���u�����t7����t������x��<SQ��¨���I�_z��tl��)M�s��?W��J��d�����ۮ���C\q����<�_���x��P��`��E�n�]��&s�2�ˤ��w��#����!a7v/��8>̘;�Ӄ�����pw4��H�&�q���x�Lt��5?�Ƽ7����+�&�A����}�&�@� �ǀ����Ht���4���5|���&�����TL�����i^�)V���TҌ()��Ͳk�{��L���>{�U�;�+{��<xr�J��^�R8��+���'bmf����9>�@�Q��SGC(�O�~����_�%Q```S3c�84M�]kF���ڍ9�S������?��3wl���SޟA/ŕ���k9as�/�����=�9 w�p�igX+������ˉv,弓�����Y�Ӥ�<6{\�(�L��4,�׾.�+���C�sL�~E�@�m�x���{z(�Ꝼ^7�o*���Ӕ����ܬ/��Bm�(���r� � 0%W�J�e6�q����uZ�}��x���1�=�t;���� ����E��t�6EOS����jT���{K5Qj� :n��2X�>W�6u��*h��6���x�~�