XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ƥ�A��|��1rD�����#&,P�q�=��H����In�S�'t�'F�D6��B4�滃ʈxe���L�N���`�Q�	�������]��\�޶�M���.�8d_��Z���e� �kM�"����˷J|��ː0	��-D��*��G���?Q�8K��{Rs#�{��P�P ����7Z�ۇ��[a�����E�IO���\��i"=�ǅ[�O�$��%8��[�3ۭh���	�+�5ϾaԴ���0~W� _[y�h�NV�n�t�$��S���t�K("���㠄�ۛ���f!��
m¥��u���L�m�HaUey�d�lP���&2��}�J���8�%d��H+ܜpu1��`��������dc�@/����yܢ�e��~]Xfq]~޽E�T����Ҥ7h��k�dT��cC:O���V8�twh�D�u�DlS����쵓����J��wtJ�Jq�A����3�O����+N������Iw�3�~'�͐����yiJ=�*�׻_��n�b�~��^���P���n:�7"��Kf�J�v�D �����+yN��8��w1U׬d�m�SD��d����*.0{�}U!m ��P̊c�~��9{+��-�:�EX��M/#�Y�Y��=���$+�Ӷy}U&�Tќ�J�,E%e�elC)յǗs&,d�t�B�bhy�j-��kb��(A�uF�b�M��BXF$��&�\^�����W=���z{��ij{J豒XlxVHYEB    1c02     a90��@!�~q�"_��@�ƲrϪ���H��2=<�kĆ��UN�cv:���z�k�\c.b��)��]�w�D��9�A㙘�P����X
F�H��9��[��C���Y�wlαA
F���`I.��G@�|��$/5'���"������S��l��E}	?�=Ji!�/��â�8��hǝ�7��	��8d��W3bK�U?{t�Dq��1���֛z��vD�q-}��F'�L����WB������텒�=$����ѫ��C���]r���x���Z���G�r���Qc�lϝ��;�mK��=S�n��_�(6�Q_���|��Ğ�rX��<S��Y�����z:W!�S��/; ����cj7�(�9�|��w���D�cᐹڨK��n������8�)��Ĩ�GM>`��s�n���O���3Y�y��*��X�!����\��UR$N���ȟ�{Qf�1�r��_�Z#N/M����$YY�_ �^JwlDE���e�Xzv��
6%ы�1�go�Ӱc՚jC���+�"}{c��Ŗ�4)P *�q�>-Ē�u��61��#��K����L�{�׊��e�>RWrl�)�=��E%��4S#��P��w�]�!1[�إ�C�:��4>��rf��"�DٛK�h�F�LX�n%�����|s���^ M�gT[).��&VL�	�L�Y8Ӭ#���z4�[��M��YdBp^(bvvu�l�tT敏��o�@�^]T8�7w�m��/x��/�������$e���2m���T~sB�v��m߬���/��[hCp��r�+I���b����E��%%~󌒄����0b��Z.%����/�5���|��?�mAD�Ʃ��8�u�u�Z�u��l�8^��*��[밺n{�'�BW��?�nD�@α!��t����'9M�wR�Jk�.��\�q�,DUv/s!re�M�ş��kX:s<+B̨�I.��Aרfٯe*�^X���6�
��վ!"��5D9Nb�O�MI�0ޞ!�7h���Ʉ9�fPæ/�����ꕸQ�ýO����G�⢿�w�M����˜/9�A����$�l��ˏ*�N��ʲ��a
��ۑ�7G�)�8��k���>K�l�k�Grym3Nv�*4�^0T�����ZC"�9�)9�j.����|�揳/d""_��L�J��K]K�����/���_�G�O��Ѝד��ܭ�Ui��3c�r��dّ�8VmŕW@������&�.4���c�I�������.�~af�[~(��T�����ַ���f����2��T 4%=D�8{`�>T+=�ql���2�t5��e��Ja�+��:��|��?�ԅ�;K����LZsq"juy�������a�6��3�g;��V�d�K��ԑ��79�!������%�ݏ���bm��.�"b�Sl�O����S����7&*c�.�}�-�X�C��:�{���y�F��2ET!�r��cތ�j���`ޯ��3��&�Aoj��6��	[C�פ���[�XQD��l�J})Z; "}�Ng,l�V^�hy��%�����*pX��B�|��gvߎ;��v�[��P;B���Q(���H�
�l��QA�ڧ��G�L����6��}��x�vĒ�_��S���to�����>����sJ���жAw���1bSIw�_�ßA�Te��
������Xp��S@�m��ѳ���i�֚qAp���]�hSh��w(u�%��W	ؕ9:ih����O�t/��<�ס�N隡������RS��G�#2���z3P�����	�P�gϢ�z �}Y���eOUz�~����lh�q7̏|`6O!�-o=C�>" �曾���>6�S2}o���rP1�?D����%��Ĳ��%��vWm����},~���K�cW���Rz/M'
�:C�"*��[~�Wq�����uX-���4����:������#*ӄ�`�P՟��?r�Â��r�0����u�5�[++�;u�D���+���I"��M'�܅��7ۮ�
�N��Z$e�je�r�e�X[\5��y%�<��H���3�V31�<��I��:!�G�t��<��FKpK�S��Ȭx�y�K��ƀ�{�~*&B�DăjYE��>�z���c5|�]�k=K�Y���dw�F���~Ps2o�	 ��Gy*����` I�HD?���d�h�c�g-_�9��F�@q9F�:b��jT�f3#�~�%��ɓd�>������^�"��W��� ���R�����F��z�#G@!pr �9�A�a �A�E=�@O���?j02��ǓV�Df�So8�r��\DȵST�/��Ö�:��(
X����i:�snw8��R���SG7�٦�vP�Ґ��,�s��Q1�V]S�;�@|�U���N��q܊��1���oV^cq`Պ�M���f�]�8��J$�Φ�K������[3�I"�}⢾-czdL��a�T�!�g0u�;���u��q8D���6+I��1<_��]?��ո�%=	��E=E	�ī�i@�5���]c�p@����BB�ҝEz��i�]��}��`Rؐ���NfH�s˨䉸���W�PW��� u	� �|-2ԣ��^h�t|"S�P�6��a�