XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����5C�(%f�T�N|Rd�㕴�~C��e_�>�c���)C��,x%F� �Ψ�Pk���+��;VU�EV�c�ǈ�	�"4��~� MQ|��n��}��E��k�a��P��ZX��0	5��Ȏ���6�����b�m��	�e�f���Y�B�ш�"���_�s8��� %n��R��|���=�۬���g�u�8�fnf�x7ʶBC4�;AJ��g6pٔV�����m ��\��g6*]yN����=`����"�<��_ ������m���<�Mr�]jvJơˎ�~��C-���@,��{�� �:�^J��%X��?�~�K@`a�/ٙ2�
"Mxil,�\̹Bό!5�"ƼT��]ݽ@p�\�zR�Q���/x�x"�:l��ٚ��kU��d��߼R�Z��܂�l뿳�#f���S�3��O�}�1��ŷI��p���P3�&/y�]����C��������U�mF�!��x�o]OTK�:uර�f���5P��&򯏵L�b����+ïaH󞸈�y����!YyNM�a�����uB��k���G��(�� ���*�jE�k���He��r�gQ8�:�5�A�V�Ⱥ�k�7Yf��V9�/�)[��b�j~�����d�9��M�zGq��]������\}��4�:�~��LޝY���؉Ɵ�����+�@I�b_� �����'fF��@^�
��n��9%۞{�(���7�J ��+*%L?M$5M�A��;=;��lƇ̻��w�'XlxVHYEB    435f     e80���?�����d�b�i�z��;A'[Jj�~<o+��@����{���m1=���ʙ��<��Œ܇u�;]�,�;�$�FXap�,�%)�Ê��-O�L�j��s�8�E��p��G� ́��E�����?��V����˳��0��{j�6|�>�5�йaVsf�t��� j#h��9X� LK��ae��ڀ�/N���P���ڌP|���E�e��@΅,�_��S>$�`�ZoEɭ[$�ތ4i�ΉF+B#��'�!г��[˒�4�r����}D�P�_g3Lm�y�W�֐$ʂ��H�&{�c|]'�.�s���0Ȉ�h�� 2��v�6���d�{�������=�;�D	�n�w�y����|t��l�\�"��i�SW���p�
^~ ��ϭb��<��-�қQmu�I5�7 q�E���c״�[\Co֣SO��f�gxZ &�8����h�9�MV`�нt\���;�9;�r��0@���x j8�v��ص(���E�%y���&�)o0J�d������������C�Q�z�Щcv$�F�w��JR��c���w
�|�\k�k2q)��x(A+H�����qk1�m���2r��Ѕ�<�G��P�n�L���Ĝ��� ���M:������FEݎdH����mN�^�)L�o���y��K�3t�?�����m���S��!Cp�?\���z�;��^�32U(.�A�
�];A0�8��� ����.˳�R*D�F-�<�����(O���"+�-�����N��s���:VnJ��٢������,L����nm�f���^ʫ��t���'�H�D���Q���Բހ���z�󞺑�g��f����n$Zt������(4��=M$�qTf���֙��;��Ӈ'g�OM@�#��m��rIc�HNDa3t ����n'�׮������^��y�17��͡�f��jqC��^��rV_��h<!�^<Mu�Lȡ���ё�������HH2�:T���C:s��9?_�S�*P�*�n	�b$8}	��Փw'�'�r�"��� ��`w�JC&@�p@�Gmo?˿�����4C�����_U��]Z�{{u-�\�u�A�����T�'��r�x�9�j�h�p�@����N�{Au�1�p��7��qy�☃_9yavTq9Lm��Q��	���g�����>�$�sO	����� �R��}���O���������cw��FѦw�@���*����z�zAG��3�c������8�{�JV��Yw���/hqg���%Q����� �ƉU�>i�[��z2�m�!�U�DT&w���~�tY"x�|�������UJ�a2vs�A�9�7ה�Y�x>�~���g��ls���3�U|�G�V���6+J PS���q�w\C��#T_��?P?v{3rK8�/�#�A�5����)���ɫ\�c����Y��<�}��}�kn[�c�)��x��M�	;��Ϙ��}����t��\s��"޺�)fX(�ͳ��9������e����rt�f[��/ޝ},�s���f���Я\�y��|F�1�������ק� �E�|�+�Q#;���ǽ�a��M�މ��Q8��,�{�������
gm�>z<��^�;)c'������T��$�#�Y����C>!������E����������`s�~\0��"=�.��bd$����+h9
}�W�6�k؍+g7f��X%��{W��5|�s�pZc���!�{QHXw��Z-��V��%�d��~q]�� ~c�M����O������k��v	��HMDdHR���=sb�ğHIM�����=he���P ��|pb�/>ۗR���C�M,L�D8��ꄈ�Z������Ւ�Kb��uAD����ӡ���o�f����M��L	�o��:�#���?P1�H���y�����ˁx��E�5t���*�/�������MQ��1���P9wb�թ8�@؍Fb�Xa��&@�w����o�#cD��S�|B�����b0�ϩ��o�K���D�#@��nZ���$�Z�+`G=��;JB�O�kk3&��2u�- � t��D�K@N���ʽl+�q w�_x���/=a�O��?VʔG� ]r}�O���_�E�"z�ki�G�F˲6�զ���~��0v�&R7P�?8��X׈}X�(��⌭%7R�(�s��р��.���:��J&b�?'�^L0>��q��}���m����PI��\�1Fe>�J`r����)힄�bN��/\D���]��e.��z)�f�t ���M4���ɓ�?H�;L5w��u�"r�c�(e����5�A�A�7
]R�{��N昗jgk9�>�$ν�� �7Y�MCD���9��w�ioh��+�����H����F����U"��l���Tj����Ú
�!8��VG��ɗo�qW3r���'�l�`6?��i�.��Gְ��ʣ��X���[����ا8�,<�j0�w�!X�&|�����^d�o,,��&����P��qض�a��%ۜ�1�Ū�pa!�k����þ"�A8W��~ñ����N�K3�fB0�*_��u��^L�f��2�L���O��]�퀡�G<��L�(�@y�8�$�AS�qd�+�\��@iM��&�ya���pS--=��s[Dp� �Ŗ�p��6#�-����p���$O[>���
ښv�ŭ�U��"�ā�QQ�fh��Z?؞��)B�����l]�$�%�Ǜ](:*t��$;G'*ޞ`��Et�����	��^����&�*;�^S�i�j�{,]Rɛ�.,;�)��Scl�2F� }��#`'�U�Q��.$���zn-�W�v3�=�n�)H�)�
?������J����혨\R%1�c�w�&�O~�?a�tȰ��*mLO�� �WU�\�9`�H'����h�{�\엧e��ŵ(���x��Ѿ�ɴ1.1	�(S�C3��[Yި
��M���8��*w��.l�7G1>3�ɶ��'�Y
�98}G��ςOU�!�d���Þ�;�o�tH�����3b����~B�A?\U�B�=�i��S;��An�O�Eށ��n�~�$��6x�ԂPu~��Y�5�=�Q�~��H��|�dJhM�f-=��"����9UY�N��ݼ���r-�<���0��x�l۹[Dg�g�|���\#���L�j�:�!�%����T����ب�J8� {"�a�g�������'��ȕ�| ��d�@��w)֖��eѶ̝�%������7�m?��.��N|�����IL��?�`C��f����50�]�B��-����8�ԕ��~�aȌ
�/�ߴ�\�����r���ésq�O������TI� [��#��[[Q�(��y�|KW����@�h�ZHҝ����l%(i�@�ElL�����f�%L�e���V�І��)��aGf{�W���b����FhD��z"�u*�q�3t뀹:La��l���;�%Xō��EsuS*rjؽ��T�X��a�ڈs�p�O�5��`�7�BT�s.�����MP�ĉ je�@;�h8�HK|FU��������6��W�I:���hG�������������s�g�e�PzJ	��xv+�