XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Z��u�T�!���������͕.�[��k��<�
l/v[Y+x��Z�8OǮ��T��_Ry��!C��{��3�u�����B!޲�Q����8s�p �����,Y.S��AD�θ�p�*)8m�!zYs`=y�N3�?`�M	[��-*�9�lv��A`"�I8٠���Vd<�k�r"���6M�'�)C^��:`
ӏ�@ڤCҳap�GvV��>ǅ I).�L�d����B85#�ڲ�[6ғR"a�|������xs_��K�~�t�[Y�Yb`����6Z;V�|��2�C�#�l^���w����w�z1/�s��2\
�'7���Ԋ�	d���S��4{(��%:��i?>=���M�'�&_�����!�)�k̠l�z��;��21_~˘SĦnk��;�T�ȭi�A���tX�9��kXTFD��#s��)��W�|�}�wV(G~�AH0�����My!؟�i�z�7��g��c&!���w�]�3�k��{����	�wN��rw�8��j]���!C�8q�cc2�2R��}��&8k�:ōA���(�G�(��j�s3�^y�j�^*Q^wُ!��'��.��������f��(�7fY��Q����Io��ײ��)�� q�U�ٺ`��`�'Z�W�p�a'��,{�pms���X@E�j��J'1��� w"~�пڂL�^�]����I�i֏|2�&N2V��|�M ј�%���Q��w�sȚn�����/����TH��XlxVHYEB    196a     8e0oh�8��\��e��}����{�'0�n�M�U��*�̓��G��!�{Q0@�.�����e1�Gؙڝ�#�=H+��gʻ��#Ƈӵ�z�|�?͝�Ig� �����Ş�n|��KAѼC`� �
�)MF�WJ�� �\�r�ο�^0unAW�ˇ�e��ƛ���k��]�3�c3�M�_7)c�5���^@R[P�(#_9",��3&b��3A]��+T�����~A�������Tf�\z��N�I�*�����t�N�`L'���R���3u���"=˙'g���8�ˑ�*�3	i��,���NZ5.�Я�b�OH�
�ɽ]��=?�c�Q�Ht�I/	bd�B�!��oDS���o���� j
C���B���y�j~�8ر!���H���~ƒ��e�S�����Q�LD��N�d�ǰ[Cv�0K-�#�	���'ek�ȟ��R�~r ����w����=F���&�<Q�_wg�-�cb��(ٸA���~�q#f�(���1%����"�X�A3&S*��"``!+X�X���)m�|�O��{�- tI� Q�j�n6C�C��&:*I��]�{ĕM�Qq�n��*`��+��/k,N�
���E& ���&pԩf��L���M |�
��_ⷈ��5r�K�CY~5��|�aT����Ǚ�I�Ʒ�ⵘ�;�]���efjJZ	�2�²2�O�"��%�X���3��^�����Fo��".Κ�*uS/ꋚ�c��I<'��1���n�m�iC�̶��4�X7?�M/3���'�M��)D4v-�����{�g��,9���cR�}7�<8�cW����`�1�f�����m3i���,m����������yܴYO@y���g-����Lk3}�ɘ��<�3���h� �Hp��d�O�'#v��"�4��em}��Ap�j�ҏtj����#=���`&�w�����Vr�������}�z�>[ގ�ե�����(l�9FN)3��-�4l�A?�A�-K!�E���)�ߞ�p��)���/W�x�nB��S � D*���Mq�by�`��S�-��΁G��A?�� �E@]S�H�S�z��'�������i�+����?՟ǃV�Gtm�Ef�F�7m5���zk�c�X���2�	��nL8OvaZA���	ͩ�a ��s�R�Z�����O��p@��HfQ�^3j��E+��䅣�?��K��H��K]J▲8�[�s�u᪹ୃ*3����gHPl�w�4#���i�$���Ѡ��c�yv�8,sl�J�Ο���EQ�}��P����~L�A��٣��(�J�2�7&�U�d>��#L%Gj(S�@�������o\��D^�����o��O�(�����+���j�Q��Aӷ���_�k�J
wF�U��1Ё�T��u�|<)��ZWo�\T�nJj0�,d�|˖`=I1�S�#��dJ��I���\�]<1u!�ۼt�x 5�h]7܈��r���!�	0��Iil8R}��R��i�0#��~L�us'���ֵ�z.���!��r3��<�_zysk�	�VIُs���@w�����;Cv2����D���	����<T���h9؟��]{��N�������(�z_H�~�bAH*�˱F���>��g���(([�3q������U�wwh�@��.����f�t_@ޛ����M���C�9�O��G���v�g���K���=sQv��t��`$��Q�Fz�x���fͳ�)�Z�νҰE��=i�����񊆛}��S�ȳA/�ܷx���Oǌ�t�#�>Hs�������(w� 䢮!�����L�{�*֠6���V�<��p&F�ڪM�6��gY��l_�a�����WF���U��cT*K����/���!̘'���C�&2��\��k4�߫�s���a��$�G,	27�sSCB,�/+��8h�����{2Mf���s�j��{��M�����&�&�|���.�d��{2\n��7f�=�:���e9�zBB���)M�jز���DU����9,�}��=�~��b�V#��Q�H������׮����}5i�2*W��nx?�=Y�'k���<r;����X"x7ʷ}����Ζ��1�nj��X���n`]��v�A�	\9S��Vpa3F#��c�x�1�Oi��@�t����]�;�Q�����_iLL��V{����;�o��z�i�Q�()��@&�ʛN���N;|4�h��