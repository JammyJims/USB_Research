XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M.B�r�O����t7���J���e���Y&��3����z謍`�S��}�N�'����R�F���}e�k�<�iکA�.cvL�'zw��N�3A=�<k�e �,��U� ɄN���p�x��5��E����w�� 0�UVsZɣ JaH����[��IZ����֧s���!�6P-,a+t��"A�oj��Γ���H$��
��ᩫǜ��Z .n�LƢ+�:�gV������C}��D8>'�<,������_�>�Ĝ$���Ӳcl���:�#.g �/�ں�[�TH��P��m����(*����;�k:89}�x���k�+��j�N�x�ly�z6x��^uw+&�/f��r�Z�B�h��:K��þ�$p���+\,���_��c�6��'l5���V#@�K�T�T���!5��E���⌽l,�ѫ�ۢ�إ����H���܊�o�Jp��k��d��N����5B�*;��h��廒8����]���9��V�̄��jS�*���	Bn�}��4�O�i>ԝΜ������\?��zA8a<�r� B%�vIܧ��OTq�W�/I$s��[:����`�p�ۡ���{�'T
GhS�wO���'N"�?��A�Ʃ�=���N�r4�(m����&�Ⱥ1MwF(仺���t}郚8����"�|���r`����i���5�$��]�ګ�Av�3_���oC,\ҹpQ��Lbw�:�c�}�E��*�~�8�7�d�pR<i'?���F��/��v�/XlxVHYEB    fa00    2800���S��Ż��&������Zx��<�+�����E[;p��(����n}�4����m�[�>𼲲iW�(�ӡohS��O�{���`�W���-����/�����r�4%�:/:�FD�3|��d�X�V��ݚk�9X�a�.�%����#B*�c�#�T��E�
�ߒDr'Y��P;���7��_@�0j7�aיW���ĵ?y]��
U
fX�'�NJg!���0�-��1]�b(�!��Г}��aX2*�h�'`��T�m_�� ����� �֕$�g�� ��	D�������:H��J�y[윩>�2�p�=Z�u<H`�ðk�+	��Y׉~c"ͫkc�3�$�8X��R���b�Րf�v�c����e}M�Aw`]��?;p��|���s�����3{8?h��<g6��Ϸ���zB�ta�W��!�Y�c˄ΩuppS��vV�D��̬�ú�7Ҽ�Y���)�|���Q�g���Y��|]iy[ɽ���
T���V�lߎpߌ&�Q|0�[l���M9����D���H��7i*�9*���!�ţR�L@1F��fU ��b��aS5�t|wj�8�����𝫈a�~L|�4w��S�w���O�vR&�1f���U+\'����0�y�K>�T����P~v��[������]�dz	�Ɣ�ғ ���Kc���j-5-�iJk �o��z��"szK��)G B2*���K�G��V���w��R�h�4���C�%lD�q�^ơ��������^a��Mr~�8�s����ī����t��k����} �a��XsS^=l��jo��,����J�Ʃ�v��O�G���!@�}>'��#��e4�w`,�g�SL��l�������)���Ⱦ� c��.���&$S����M^�����.S��Cg������jg����2��B�j��O���p��$t��<�^��fk(&?HJ�p{>U��@��K��m��0���3�
i�iZ�w�8��i��0���d&:��ٕ��� f�  D��Z6u�W��@-�?h���FT�W9%΂_�������;%���U/���1&�Y�r�`VƉ�S����en%ө l����"�\q�(E��$g6��{��>�4u�S��u7S�������FC��U?��μ��P���9"?�E(�T�Ul�ѹ q��=J��Ė�(����]v��8�+d�ͥ���=1�ʇ���']/b���;�Z���W��+#�k�k�(CD������~��q�:�@w���a�^�����D=&6��~����"�>����{FO�/���1Ť��/����c^o�C��C|��*+����I�L(��Dh�̬GĠ���a?�9:9�#/ya�;�N� :��Rj	�|XZ�N��?�ή�h(�V\�7��Tq\m�LZ�ٸ��5%X�Փ���2��i �m�� �>��d����~�tg@�2Y��H���#XQ�g�6��;��&S�1tƬ+��n�H�Y�1��⻎���R�{����]ԇ7����5:����$6���Fy}�;P�91�%��R�_i��p��ׅ�8�uOI��P��.^r�o�x�l�R��b��pH�v[���@G��h�rgm�M�6H�����kGQE��3.H� �J���t�Ӷ@��-w(�Ђ6~Pa��r���	+��2�$�r4�荎����S'���]Bjq�����o06\�7��{4��KM�,�qB���}�z�����]��p�CB�R�f���Ae�
01������ -�'Ĩ���N�]F�V��O3�^��"{WX3RI4�.u�a�α��A*�Ȭ-�NI�\kڲ^.�hpd�ӟm�<Q��^�%Q ��@b7i5(����K�ۂ6��v��w�e��j����B��%��t�)y��B��;����A�Z�&$��[<�j�;�󡗂��� �Һ�{1*�o��Ҝᗿ�w�~���,Г5�3y���H��	��
 �	�$�m߹��JH��5NLnw�eP(�9mgqn�B�OM$0��|�V��
�����<P���������%��$��Q/
�0̔g���9˔*��2q���^S9�y?O�HzN��w�<�q�{a�DU�y�X.WB������;�A����]����a
����gv�*�s͉�w��W�e�75(������H�����^
��ߏ1i��>����+��!N��BaAG4����y�Pԍ�0��g_�{n-�^�G/�-%X��-%��3F] vsz4p`���}Q�LZܾ�붟q�#�&j���E�5�h�>d��4���kR���+U�Ѐ��#)��a�nC��}�)moں�7[�W�D/��M�AM9�je�#��F.mC��0�.,��2���k���nI�t�����12r�@ U�@A��֮z�nY��d�� ��(�R�ηe�\�y�ϖ2ǈS�!=?���������d��Ց�,��D�`:⴫= NC�t �Gh�� �u&��aZ� ���OUԟ&z�\��K+L�|�Kq*�g�f��\r�m		�x��K�ŉ�����od���#P������J��VKr����x�g��(��}~�s"o���S����j'ګ�� s?4D�1,6Ǫ�/D�*���Xe�k��8t���zs�	�<�]���f���[+�1mc��9�`"!&�a�/h��I��ǶJ���u��\;r�^���x�e�i�X���)Oo��}�����e��ĺ+v��oF���_��E_ۙ/*����e&��d�ܶ*��N���S#�9�#\��Ni���M��t����L �L��Cg�h�_���jU�f"�ıIy�<+����q���/~���o��B><8�)]@��j`�������O*�KگG�tSw<��q�8'gd�RݻL�9���&���K��3�`��v�1`�����(��A5w�G%������gg*�DEEU�a}���D�>�=y�YL֫/��T��I�9H:�M�����i,����>�jpJ3�[>�T�e��(����YЦ�.����0��f�����`Va����^*ɶWړJAr,���;NMr�RZգ��$ ��¦�(��l�n���^]1�~���ʝ��<N�D�^���ws�ȒYV�&fgK�U��W��L�N�֤�l���:P��.4S���T�6�x�=�+��F�O��U�Y�"��LF!���*��-}H��y ;�D&�����i��=�6ܷ{[�U�K�ur���.�A&���}(��B�~j�đ�A�ID�%�l7ҢTs>��-Q���|M�f���l�r���ũ�A���oR�'j�.^��K'��C�ɢ�&`�J���±Пƅ���[��	eK����`J��u�4k�*�O�j~1�-�0��_��d�,+��Mwnk�'�'
7��#yGN���H�����(�Ǝ&�I�O �d#Z�?4n Y?�Դ������|�w�;�ϱ�S�B�7^M
Ѱ7Z�!��
ܪ��aÈ�����&��=��ed��B���bն(Vk���g���2΂��EN(\��Yo���%�Z7�޲Y!L��%M��Ǎ,�P�b�����p0�����_\	6yŲ�L�9�����ɬ��П/���`\]��:���צkش��m(�\�����C�L�nB�<��2x|���ϣ��?�4�ف��YYv�' �QXY�\oV�+�Lb�s{��+{��7��q?�tEr�,���(y!p�,���@����0A��z��C�VU�c]�~X�Ӹ���9��`P�CfJ�ક6D�_��IR�'�����C�(Gd`ͱ3V%�7��b}��п�R��g��ͫf"���+�Ϭ��@��K� ,�u'���Ƙ�Os$�9{����n��%���h�����:#���6C!�t����[ح$Ź4W�a��Ln&��{�1S�3 �9�|��*J�	����Ueʋ�GŤ1lxR��ƨ�7��-��,4E���s�6T��*�z�E>C�s�8�[��py��@��Aķ$o&y3Z�%r[��[{��e��J�w�����L�ؒ��ھ3)��C�~���O
�uJ�$���Ġ6q	��P��]�tV'�,Ƭ�0�)*�2����hU� 겁Xz���1��qB�4�sڞ�V���9�}� }zm�%�RGZ�T���7�.b6�v$�l��`S�S��6�FM���&G��J�e��aUl��L��9��# á��x��|哵l�-;�L|�~�m�mK4ب2#��V�n�\Pp`T��U0�{�7Tl��L�ȋ-�T�`�����C�(@���E��JC:�=�D��� �Sk�D���)�d�~j_�l�K��?�#���e�����(�t���?^`��S��27$��P]wU~sagN8�$�>?�������o�O,l <�,��E*b(�K����X�+QY9% �)z�(I�WAs;�Ր���!)M6�3t&Ny�Ϲ���8���g\����6�2c���X}з�I7�!�wа�j^{���.6��"xncb�WMq-���ЀW
䋁`���n��)���0�j�˃�a��z�;�:[���D������P�_����2�H��S��r_a�@Xu�$�=<�X��ؑ�M��?
�=��H���BV0�����m�k�.4ls��~5^P�՚vdk|zD��\\�]R�zV�����U�dq|��I_��)�<Ɓs����1�q��"5iL~�_!J z���/����t|T�Ho��t��o��@��Q��g ���h�U�����?�M ϡ��������[Ԁ>|��s{&x.(l��`&K��G�D�.��X����o�����A��Y����ʕ�������dC�N���	�!P���a�W�˷Wz�z�2��g#���� =�Y۝�@���|Htbr|����a����]6��8��,1/�C��3}�}�wm��(��|���/��:�B�7�E�Zf��=$q� t)nw�Ki���_1�
lC�R�}Q�-�6��ܔ6H}1רD��)l�qR��|�<�Eo���^6101�!�P�R�޺�z�Z���	r���|�1ΓL��T���j�K�F�	�u��v�����˳����$&��;�mdz�pU��t�+Re�hG�]�"�>�OPW�/�abW=0��#�פּ.u�fo\'��i{;B��y'��zD��- w�Y�{�	`�*��e[ @� @�.1jO�����3������ ��l�ƲQ�7"K-3��lVt�}�;�`�T=�[�K�����A�P��C0��K�ܝ�М[�2��E��J{�F����o�����R��M�q�Z��*�Mq��p��ms��*�4�޸��� s�SV������~�4J��Q�A5�Z ��q25�ޛp\=ٝ�����F�=�x����_w�l�8�
��uu��	��h2�:����}�L�̳�,����J�!3:����6(= V�g�%��jym�+������C�d�uZ� ����.���K��R����8+�n��`����&��������'�.LA/y�$��u`���n��Eɞ{���z�� CnC$�j�����m�D��^� ����LG\�:`T��9�$*�{>��5찚�����$���:�v���v��P��ֱK��R��ѿ[��k�?[�e��Մw�Exع(���~/+5�`x��4�������Spkr�S��h+�Գ*�Ϛ/>����7�{��I�6U�騞�B��$�������%'{ux�f6z�s�]�Uȝ��.�Dԭ~|y �h	�/o�ƍ�5fl��B�P��e���J��߻��K�4E�qo:����\�����|T,fR���bBy�v?h����9�������Җ^/U�~6mC��z�G��]�@�*<=���m;��B�jL�����ȝ��nuH�3$w?e$ʨ�"fK���3��K��pZ!M6R����{� ^��aR��*N��	L '�����.ޣ�8זN����34��W8����%������3��f��Ѐ*��*�i�s�f���O3��_F�=���1Ps\�:�H�:���c�,�B�V��� ����яIkI���q�9����|S�zi�5�wW�"��O���C?�D��#��"]S�Ļ�U�X4���.�.�1���#w�c�p{=��q��0�/�D�E�5�,��:��r������|���@!���yp��N$n!��s���r*�Ԩ4����(��'�z�Tq  J^�$�a�����^��qL�$�B�_��Ѕ�,&F��e���eh��JÛ��Q%�KY���ۂRE�6��^�H]J}���wb���I �n�
��Wb(VDY&���멠
��U���|0�f�C�z�%^W�n��k%�#>�tF�vN��.�"[=��QT Y�R2���\�57$�i~/9P�nb�o�&����2ʅN�''���^Q�5�01�����j��'� .��A"��G���g�c[���~��/Dd�T�/���4�*^����ƉHs�8����
��y��?J$@�Ĳ� �C�X�Yt�"�ew��q}�jq�y����{��'b�Q�slZ?X�(�M	A-��\
'���8>V��UG�������S�:C��0��L}j�m�H�^\�lP��<'�kr?��P��>g(��p���O6��G����y�R�g��_��ݛK��_ah<9� �"Ǯm�l�,�_qER+_c@�N?�忦�һ�+��V�<��\��w�_o�z}����&�`���o¦D�;�f*dIl!����F9&Bz���Ɯr-�h�y��9ô��bD| ^����]�؊I2F�%V{�\�.Z�Y��`%ugk�R�+�+�k'R� e2b����y>�� �T�Le�e��M3=Ұ䫫u�!�~�k�0�� ���)��e �r�.v���[�����#(8��E�A�S��zq�70��\(����|��g*�)��3�{�f<Ѩߧ?f��u��N�fG��/[fw����"�(����� +�L�VsX����d[@���ʸo�y�=)�t�z���qF�-�4j9!O���~-lP׿�����m���yw�;�;��/%��]D<���}�b�iypӟ�<��K��c#ŏ���z՜�Jɠ�z<7&ПR�ɼ����4��V�Q�iHY�7�V䚧��Ng�n'<R3F�|��=�~BA��Tԇ}��4��I���pąE�2���]��[�y=���-��o�ŉo���$��7�3����N}b>8gHk]�i%��`��6V<g�]꩒�WP!X�Z�.�4`g���X��mD�r#"y�|VlJ]r��ґM~�6�8����(�O�H.�r�Ծ���n=}�و-�g�D�t J5��6d�ɚ{��;��b�0�4~'��=��~.7���oU���Z�"�cL�齃�8��Ƕ�=q�}��űW[�Ӟ�F�p�&��L���8�`�oFZl2�}�.��GC�N;}�|h��U������\5�f
dׁ�9�0+�QPR�GBn��	��8��N�S{b�I�
�Yh�#��,��.��E��'=I4g�D����V�gC��P�*ǃ��\� +���5¬׉�AP}ȳ�|��#	�b!:-N:��}��]e;��@tC:�I�129��M��M�>\��ڌ��Y�0�8]uN�8n��(l��>oO��%IX4��J�㘈M���$M��,���;� a��e<�]��m�
�R�����y:�m��'J;��y�0��+_�E�z<h~����tB��Cu�[q=O��om�_��l����Ӹ��{)O&��o�l �}�Y��o��;7���>{���ic��+��Շg!̩��-��1�]�o�ݰH�4w�V�:]���Ԑ)lYw��O�p~��daDEN�!�#�9ףh%+�,����[�0:�xN���&)��I�0?�-5��I��2tIPu�"N_���՘��ʗ�����M<ّ
����l4s�%y����s��S���.���(}A���N�R�"�:��URj���-�M���u�;�l(^���Pq��'TW_|�E=ǰ�/��Z�Oޓ��Ip���;���q�����4c. L"����M8S����v۫�Ԗ��� �1��hH�_�'��2�R�I\_����Rő^��G-2J�����	MFr���"Eȷ�]f�i�X�=u�����m����9��#�D�����Ť(��٫V�Qq-+I�Fw�*_���vkE4`�f�\Z�~eMȴ���i˞zB��E4\A��6�_֨W�|C��Z�W/��F+tZ���~<������ǎa����E��F��C��&8b���k�?,Ⴭ=����(�Iq�@\�c�܁�ʷ�b��ze�ڧ�)"�L �Gܖg�<4����Svc��?8WV�R���1�Ntx�Z�V��iO��R�����*$��j4��fj!��1-�����g[��uT���f��?��@����H�����@xU���=Zp#�sŅ��{�/�i��v�g�9/���@p�>��d��c�t�8�%����HXQ�z���ʪ�50ś��ߔs�ҽ��6]!�/1�5�T�`"AK�b	�>pQmrv�f�s�0�_ܚF&F��q���(?�2��3�g=R�!KVx-�	f=' \\�������
ՠS�f�YN>ݥ���a�®G*};i���$���!N��(h  .������-Eo�k�3o+��Q�7���}"�]�lO���̓x��/4�9Ş���摺�͕-U�CPw���W�%���y]�Z�6ȅ�Eo�+I�C��b2�%���f��k7a��l[m�C8�"�иS�$q��ibկ��`/�"+�=�/5^%I>S��ቌ �@�y^���PVS���=��ZG�b�tG��Ni6�v�Ժ�Ş�wDm���,�������%�ܘ6/K�s+���x�g�Tx���������'��Yy�����1o)#;k�)�4��%`����"Ύ$���i{t"Oa.4F��>���O�ΰ#l&��p��-z�oqR�=��s�_�^�J�W΅X�n��6�-��(Xڥ��^��m�һ$Mv��.�#�,��������4%?���/Nj`�b1��9��UB��I��l5-e`&xZ���M�S��9�%��d�#��
�Ma��=%,��&��q6�>#��%��v��b?�b2��j}���5�9��_%�IflU�D��u�/-pv����yK|q)��C�C7�Ҍ,����ZN{�C��!Z΁��z�>D���k�AF`5Zs/�|�tS��2��#9/hh�9��w6m�$��ԷbӵDRN)nDa�9�Lz=3�/8`�4�Y_o�d�F�ى��{�[`���#�L�����`�o�z�FS�}��1k�KLQ���l��M���J	�3c��R+A4�=+�&�Q^vs8y�)�Ӄ�,Q&�#��F���I�Xߊ#�	�����s7�Ơ�)@x�:��^�9�_{O��\-d|��f� ����}�z��&���8<*?��{m�b��߸���ã3�N���%�1�F�辝#�m���
�TL���Ǣ�QG���w�T��L��k��U�|���/¶v����>�}\u���S���M����R �̿�k@gO`H�aԡo��zl����Zb4Jõ�]�T�&b�۽e~�uYW{d�޾�\�.�M�r�;FIjer��U�d������Þ������=���%y't8�a�Ӣ�p��ҽ��	Ҝ����P�f���J�,�>n�1Q�]'x�]�y��Ř%���͛�S0��Q��"2�2�C�a�V�Pt1�L}J]�bS0�f����m�=2��~~��w����ɓP��(�"���2�M`�?��j+�,֬�L���v�8��W����Y��8�f�	��En?-U_b� B+�������%��#L�B*Y%iQ�pnÊy˱�?lw�	��XlxVHYEB    5ef5     b50��3Q�h�u����TD��"��A��'�X����-�Sd���s�5O3I��kbFǇ���;dP~D�vbK���K����&.�IK	C��j�4�|M�sצ`�Ώw��/񩫗�5Q��=�����t�:��N,�za�n�� ���v���2Ţ%x� � 6ƕ�i�-0eP)�E��Ih~����b�[�#�#����f|�\���kԟ�6pN��kS�T{>���|nO�m�p����'��29J�,u$�$��Ǆ��6�G�m=yE�rQ"hKs�-pm�IN�Rd�l�t���A���kg��&	`��xf�JtJ$�6��FH�p,����̍5g�Ƒ*nH�E���`�Ŏ&�{G�7�D�D��ֻ	�I6Q�$�l+$>�#ܟ"�Q|����zP��:��vH5�3\F����u�/�� ����J"TG��z�5��UO����(7�w�Z-��/����%�'�B^�rθ�l����5s����p26�q���ET�Τ�����F��{�B>����J!�Y����}&�5|Q����"�U ��L��ɩ������G`�.�6��\�(S��!��]`ج�k
�x�&6P���Y���7a,��aw��)f����N���l��y!}�'���B�c�W��F���n��h�}�"���Mɏ�"UgJ@0����yp���+J�K����/ѵA���p<1\Ds�gv�`$ޥ��EL�
���A��Pa�GX�<I��3ڽ/:l�f;�RZ�ea��+?�ɵxz��<��������9�!�� ���u����0*B4�K�����C�$������4����,��6���[�9�6���q����/&k6UT��e��>��xzֹ�NZ��ž��ol�tA�n:̻Of�1;.�H�F���e�x[	9�6�1y ���iB~�\����p��(}�mT��Z�\���}ȳkGe�h�q��V�1]q5i���"�r\�u�혂��Z�L�kUo��yU�pR��d���+�N�G���6����fn*�6_Ґճ!j�|k�m������i,dUߍ�F���:ҫgnd�>`��r�(����3�z�� cܶ'DI���2�׫����Su�fT��4��^M���g�~�.�ԅ�R'�`�7e�m��fgp��4��KR>�O:2��w9�{2恣1h�V�9N",V|�Ԍy�kd;�j�X�+��Q<���5�M�b�N�OD��63�+A5���;�^��Q��M���t�h��k�Y8~{TW&<F"�-�Fh� �_��S�� ����Qӆ/iSN�#u�����Ut�oR��p��W~����̀
y$`�t����[p<#�@��;"r�~�9��ޯ�O �2ʐ$�PXһ/H��q��Li�,ݔ��TY�?��/u�HK�4��IQX�l�&̻����tf�GDe����8��FY5s@ �57�+��~܏�=���\�H���ƣ��-̹��u1���%�/"���A�_�t�I�	�a��;�P�G&�ߍ�R\UQ�Jl���aU�ᒾ���c��
]�|��ґ�3���޷U��m���9,�;$�:%[S6�)_��rK�NÏO�j�H�~��j��x�O	�<ַ=�ں�i+�v2
�hĮ�Ɣn���Ź.pX�C^ �"V�����*�+�oe$�m��"������`��7gF�q{D���5�Z�n;v*�2�]h�!� |��a����`{�E�~�yB��B��E�&;H�?z�ϼ��۪ȝNEQ��ާ���?Zs��J��מl}�P/��(�R�ӑE�S�uI�ٖ�G�\r
��_8�O���9�_9��@1Is��#9��A�R6mP=)�cz�p���ě=����A.`��_�BGD�ݓ�|�<�K�"M�FM_�P0�D�B�x�lԏ��+�����Z!v�&���	��89��>�̜��>M���+����;�y*	FG�B���q>��e�>�`J�����_	��*C�.%����	°����F3򸦭ӂ~/���
EMZ�O�יzC�e���#)��c:��������*LcgNq��l���{�zy��j��gHV�ޣr���7N�uYwۖ估$z��~X D����������H�!u�RU��li�h�uKm\��mf��	�iW���x�H���k�I_�e�O�-n$���r�ƅ���2��ѣ�]`;�{R)ؾ���S�`�-y]�Բ������EՇs5 �̎�8��+W�Z�dJ���n��a��TҺ���6���.�:9�h�0�)T9�:n����r2�LA��X|+o�r]D߫�8Z�׼	�� ��Z�r������Sv$<�����+��շ��@O �:��K0��"b?}�E��fpE�61�ˈ4�W
|�=�*?J:�pq7x/�f�C0������S�����d�w��u��sH��PQ\�]{�9Ӻ�����N�[D��eBSDm|�U���g�~W84Y
��ׂY��nl����bI+�&�h�g>���5XVp�W���H��"��Ua^m�HCѸXR��Jg{؋��xeM�%݈�:|7HQ-�5�+{ �SqS��4d��|/@�kD���b��4o)�q�ft0��v�A;@BB�O���C���]Dp/�?���TB���cMsJ'6�u}t���ƕ�z&uO?���R�"S�>1A��dw8�����N��D��Hl�߆��$Gl�Yp� �qx��{Cvcht�L���u!.N���z[1�jN�vz>Cٯj�[�S����w�M��$��@�m%�_��x◮ˢ�٦N���]���IS�