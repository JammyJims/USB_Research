XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������u��},���g D�V%2rT�ql2w.�hU�D�ŗ� �Z�hMS��?~ZΘ���e���'<f2��/��Dlru�h��|�,jk�LO�D�q������������(,���y�^,��=T�h�)b_L��MF��4s9;^1O ;L��ي-�q���������+�\���ڙ�Zd��T�3s�qRa�9֍��l~f>;�߳0����L]�"�l�W:0�$_-��%g����i�w�dO����׊4ғ���b���P�'��ǐCX��}4�z��d¦��<E����1�AكF�A/![Q��%���S�;�7e��Ex��mD0����ˊIv�YD��?��!%��{����o'-�G:."�������rr���)o����2�k<C�� 7���v5{$ȅ]��HԊB�K/�`h��<Wc�UBie�񘕎��B)t�n�ߕ���{S�˄6�g����*�ӻզ�K����1&�[��1��,����cX�u_��d�U"�46xm�3� �n��ۖ���Zl��'��r8W���?�yؓ�%��7���a%�����ɳǻYv�G;3�SFDe�Gk�g?�%�{���꣭U!�5CCn�$b�{24;�_c��j�(|��&R��S���8�98z�E��4�&��Ia��a�����F�;η��<��AT���6�3�Xe4�8����]*;u��.�p��*�H�`a�Ж+��:3���ɴn4w(K�n������ͱ��#�=<XlxVHYEB    3f51    11d0��/\�
Sֺ�c,$�RWB�bCx0����'��''Y:��_��,Cz5�;����GI)���b/��G�Pq�i�+�NS	w0&t��};�j�;�c�k-F�Z��o��YK��hע,��w�0ª�����&μ(qd�ەw0��[��$���&)��l�ܗ�u&^ J~�eP$��VW��D�N���/j��*��#���K"97��h�9���}G�<� �y��B��K�P���G�3Gŗ�����q�{9E`/�����8�']2��2�����c[� 澖�����z��f������0��R���V���"�����K�:uU�y��h��~H�, L*�P��%x��Q}��ܝ���Xx��KDom�K�e��U�B�4l���(����S�Ac�I�R������O�
!yE��o;��8x�M׳�ak�*�%��C��t��R�3+a:7&�~)�	��c��#�N]�E�.u�l ��(��{H�q�����s�q
�$�W0ޚ��rS(�U�˥K �eO�O��1Z�Eӏ����~�k O߽ʰ�8]R�R[ / �_3��^�ɩ�P��Wf��癥��)�xϪ��`�`�ub�&��Ū��:�P�0����fI�����$�Hq8��h����-�ƀ5b7#���0ԃ��@���Ce�G�����r����>�����~r3i�,֙��R'����6; �%�<(������sL�lOɓ��U��E���5oF��GW�a��4���o�o�2M>�%v��b�O6��Za�O�OE���h�WL�6掣?�v��]���
���x)2�a}��Qw~��ކhPJ'@�W��iY��Pm"�ƺتW�����E���O��!�q��X���e����/���;�f�\P�ە:�� ���n9�{�m'Pgp�+�/�j�?�i��>�7E�=�m�~�p>
���K�W5�IG�T#I.�� )Z夃~-�n3TŌ֍��>��X{�	�.�:{��6����1>���w������.�F�=���ⴕ��39��g#��⌀�5��X�6�,f��(����$��8��N.
���/f��޾���Rf<���~V)Y��+:0RH�s#�@�zwܑ� ؚ��;��S�p�KP�b�a��Ǫ ���Yߖ2�J��dTى�l�{IO����i��XAs���N<Hn�0�Uv�.{5h~x㞤�w�Պ����
�i�zH�9�~SCpk�g�.��"���_8t�$Fs<�T��lϏ���s�f�b�"ŉ!+��l��/�-�¢2{d���Eʬ*.ɚG꙽���|.��xW� �]��|G���4�B�_w��|>&��B�,��x>V���
M	��x������?X+%�'U�%L�!�CR��:j�(5}�r ��A�����@+=��M���-�C���xg��$)~��87]��zS���Ɩ�27�#�/@7Ų���.��`��3R+b&���t����+���e'�_�9 �|�����nt�����Q��vH�^F�X��r��2).b.�j�9�8��7��]��z�Y;zk���'���1����>\"���3>��!�t8���o���8h�Rr��]�̣�]�
5���Hu,�,c?:�������}�G�]�ec���B>k���FxO�~�T����E�̶���kol��`� u�l�[��`������1i���4��y�KHZ/
��̑Ͼ�cYS����c�j|V-��nQ����I�H7�C�|�9��I �i�\4ahᡢ�h�K�]zW]7��̳��u�J!9��(Ḗ8�X�doV��P�7S���Hk��}	���rA��I}��Ø��H	�w�g�0�{?ԛ���`z �C�,.�������aϮ������[�6�푞d�S9]
,.���N�Q�J�U����Ӻ���?��`O&���#���U1P@t�s��x�I�M�����g���u-�/���I��ia���-O�Q�}ԀK(�x���(08���U��ϑ7j���t6U��a9i-��,6q\���e�̰x�x����К���p��0p+\��ɐ�F3��
<#kR��
�)*����.�h
'��-��
EC��QgP?�����4t.�Ǒ�k`m�×�I�8H_j�p���/�]#!)O+ Q
��o��b9>2�.�����RLʧ����%�f�k���_φ� �����"�x�y�WY.� �'b��|�Շ�m��i���o���0 �B��n��#���j� B��S�Jx��u\(���i������9/-���J�%u������C
���ec�A��]��r�m�8��o���q�
�����味Z�4~ �������`Qծ�ʫg�j�1=\����X����-]O�s`W K�J�F=�1�GT���p�L*�8["��R�4�g��ܞ��e��26�h%�x�T�% � U�	Q�m���8��5��Y\��}2ʺ׫��� w��d���������WnO$9�^�=�_�3����8�"pg�%-b���\U�c��0�Li�>�_Iܥ⺴Z�}1S��Q?����!��ONz�+��3&R�l0Q5�T+�H��_�=�ڥp�5�����i�2�����8!�&���O��퉛��}��}�q��W�� ݍ���tcg*y�*�VG#'��H�}M�a�����i��^��� *챨�,���8n����T�:FLmj_iЂà�ó�^��l"������3����s�9d�q�]dJ�%c�SYF#���z@��o����4��YK��'-�-b�g�X��^�'��6�S�tB2w��h����i����D���]P��b�%�#�-OP�� �'��p����JL�Nȁ�b�W�n��:�4�3�]i�	T�9vd(�b�W��m/�7��r�d�:�e�lΦF�o�P��@����B���~�Ll3�E��0�7�e�WN���
�o���ù#�M|��$��:��W�s�,˂E���1� B���y�U-k���]�ˢ����'9��;^�W����W��]��n���	���R�};��xTL�O�) ^��	��LD:.&DF&y��GP��~���|Z�*�WFOk�-)���ok�/o���Jg�m�h��{g�* �Kԯ����GIv:���3nĘV���X�J�/a�<茬Z��G��@��G\U�� o��Jm�˪�s�{��(:H	�P9��s��qfB����L��尻�W���1���	���G��H�w�D�$�4E�dv)�jc�[�~@{9�iS����X���q��Q�@���[�@��`[h�&��b��{-��|��ѿ7�R~���1�-��!���a�$�u�ժo�Pt	pf-�����O��V��<<����X/�Pp��̔V�D��Q殷�
��us,{ɸ�	�ç�)���-@N�� �A-P��y���#� u�I�>�4�0�?������~m̴�:�v�C����i����f����v�~"9�Fo_�/��[�c�$P�����kGw��ң���@JʎY �ҫ|�\��%D�}��d�+K~�>���[|PeYȇ�Q+x�V�h)B�% 53���16t�M��!�=���em�vh
�t?l١�=|������I�����v�b;�B�	�%NN����� �x��s5��X�r�G��S�x�i<�麚fw��}��o�ΰ�T��F*�RC�;>�����
�{��Q?�D���7H�H0�3��l���2�_���Aɧl�DR�d�bIG���<�L�)�y�Ehj��(�k%QD!+� �N�ި��
[�6*65��у�sG�*<H�	$e;Z�*��,��&$HRMuaF2�H��P�dO]xSu�R�����G��Q�&�����>���Yy�:��<@��@�JR����-��������,�Lk�[G���ӌ��zL���%s�:����7��T�g����<0��B�ė�H_�uՂ�o���d�&yÒ���Jt��J&��+$���3|dMq�����߅�t�_�-G�'�/���7"1=Rkٖd<��E�)�Vc� �E<S��rD��*�����7�]�L
|�GR.�wg�'dF�J[�t��GS�B,�2?����y�xqioDN4,O���[O�����%o���8,hwd�F���w�����qf���&D�d�yη�>��j�����zs�3��2�4�x\]�100a �K�n��*o1�8\���m�hC��~+�O0��t��z;E�g�Ni�2�����4�?�,\�Q�:��Q����찴�����UA3k��J�Ke~����-j��WG<�C�F�����~խ���]�%L�%[:��;Q��.{?b_Ì0����ÍT���W��-�*�s�WW�x��s����q���SJ�i����#Z���oY�r�[�=;���� �G�Bw�yiI~��͙)�ŔH���AD��d