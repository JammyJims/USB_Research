XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J4��WT�r&�9*�f ���A�5,+�gW����	��;�E��O�]C6�5��B�W�׹D��&������.���Em�.�\Z�o�5W�d����1�-�HTꫯ��yo� b/l��3���b�b�¦m��9������f��=
0�
�Q���$pn���1(t�$87���G�.���kCƿL��2N%?�]�]��DљO���d�T���;4h�
����g��pe,�c@*w�x $򳩼n'L��\e�1_�=�E\�H�xg@�퐠#ռfޙ��h�0r��Zb�;����ġ�ξ�T��"�l$�,=[]����>��F������N��6nu�K�f��FI�4:��.��w7�9&�b���T���CQ��&�����u�V@� ��-6�)��8 Y��+�GOOс?!+_`�����k�?*n����Ca_���'1%��a�>Hj���-�"!�����E �={\%6 �fbO��0fZ������i�"\w������giy�+���Z�6݂�oZA�F��TrQ8K>�E�B�Tn�2H�pC&���x��� �.ʔ��5��tC�܌�<�˾�Im0���4�	�9��0g��΀��]j!G*Oױ*NԐ<	sp�ʺ8ތA��eQ4.�y�s�W͊]� � ���nt��ؾŻA&x��5	��
�匊KsD q�AH����^3iH�?�>���)�2�.��U���D_�A�Q� �Q�+�z��)�lXlxVHYEB    fa00    25c0�[��>m]��
�x�=k��M�T3�ZS�,��hC�=2�HJFr��8K�E#�[g���7Y��)>�dtM��:Y�t��u �~!�+!e$8_�����v]4���oTk�OF�*d=�;����|6��'�A.Rȏǣ��Ў��:�X�gט��z�Ώ�\�>z��Y9Y⣊���?�kY�p�V�hw+�҇;�a���\��]�!]���}B��^��&xY���g%p��=�q�u~�l�+u��2AI��j������XQf] �ܣ�w�l�R=ݏ:y���5���&�+�aC�x87'h����)7p�	1?�H��7\;�m�͕=��c>��+���e�������GnG��Ss�;�c�i@x���
�{[zqe�T����E���ţ�@�'�<���jI��uί=��!�V#r�� `<�v=e�����D��"J�؋!�ƤE[`����*��w��c�c�0���'���u�5��2�5��/3�ܮ��]�Z  ���^:2w�#@�MS�{c5��+�P����8R����B$E��� ��хQ%�T��b�w^�+�S_}	P�e�g��a���)
\p����%��p�R�_9�o	c���ҴC��G;}���V�s_��gk��w�#���i#X���JT�:�V�VΆ֝9�W���'\�wdƁ�B�
�1�]RA���{c�;|q�s�Rns`�u�������%��x�5/�hP<��I1��82�"��x���:'�n{��0��\����\�SX?��X0!�w3�6�Uq�W6�& ��*e��v�^p��v�����@�U�Ru���u����2�'�#ly5��N%��O��]s�������i:+���c%��Bq=��D�;A��,�p����[�o�v��{J<�pLR���D�2�� � _О��7�Էd��Lf��-�>c�3R9����d���0����k�U.(·|6��.s���X$<�ץs|[	�HcWI��K�x#|xQ5턱l��n�Ua��uǰ��gjxE.`ڦ_=>���(KP�8ل0�O�J�b�l��]����̩9�Y-��Iޡ_<�~|ľ�K8�l�^���)A\��o��JӢx�D���i]I�oo]?�N�5���S�,Y���OQ)��}?b�B�}�Y�y�8.R� S���TxK�g��r�����
M"R؜3@ȟa8O#9X��qz���z`[;%�ݣ���͵�� ��N ��CAA�u)��k��$��������1�:���7
y��EIW�J��/箰��o�kJR,��JD�E����<����t1�r��������#� eÂ�DW41p�OI�-�Uw�,�P[�i�vq}҃M�k,�7}�^���:�-�<Yg��dvS�l�ϻ�u<���MKC彿:����ػr������;�*�9؛hc�6��%p|fΡ�[���n�A��:�����^A�$!�z?Qk�8�2�|6�2ܼ܀^8.8>�	|nN�ǤF�}|`>�;���+{�d�˾w�*���=
J����Y��c�n8�n�j�c��~[�yۿ��.��Y3����o{��n��5[�X������M8L��1��,=�Y������"R�P���8�gz��q�y��
��|�î�,�
��e��O<�)ڃ�w^�s�SH]?�v?��"@�?9;��U.ػy^�7�J���7)a�8���ֈ�|y?,t6����ŀ`V�:�_�����ms�+Tb2%D�����8m x��i�6�tT2�;c����EQj��ūYe�
ea)-�S9dQ<�����"�lq����oI�fF��;���Ľ����z�,�8�������Fl]�
4����@"�%J�\.�c�a��.a!�ӰW{���c�rZkTyP>�bߎǥ
-v�r"m4�BBl�p##i�N��u�WDm蹷��( �#�p�|�=����fQ"��I��#�'۽��D��M��Y��<A�B�eg�.�06��FRZ:�=���%���Gj�v�2��ڟ��5��X���G�X�]�����޴������F����}h���J���T��s%4K���n���2�p�war-��Y���q�S&�R"�1 ��A_IOP��a�x���Ѩ�{�g�/p�F��O@Ĭp�m�G��Vn��=�/��ׂ覆sϩ9O;�@oj�slE�)b~���S�V��Q�P��Żƛ�k4�y���0l�����,�I#�ܬ����i�`z:�����U�}o^�L��������9��6P֨S�WE[�ǣ3���q� �EL���7(��$�&�#�U
���Ӎ��W)��80i�~	��!%�p�x�ls�\[�yNq��L9K����&�*���`�����b�T��ۖ�8h��K�`!z.]Nl��=���s��<(����Ow��u�U�3"�8�����4�&u���펈���'p	;n^s;�vl�`�';�a�/��-�����齭T��%���0P�氲�YQ+Z�����ϺV��K���$}���{wz���0i�)$�H���B��+~�w,�����S�0p�p��V�ņ6����̑���
���P����Ey�H�K��8S��� �y�B� ��R���s����k�
�݀��(��h�֧l�Pn��R�;�h�t�ã����i���JD�XƨQ��Y^-��_�a�4i�}ja!6u�*�/����l)�Q��h����?�7�u�E�����dR��V�l���/NP����phi$Z=�r��g�
r�IYlcN�۞9�<���^��gF�� [�߽�cF������7T�OmĴ>�W��sY6ݑ:c�EL��:�p��� �J�t4�b�0΍'-�J�n0i:��{-p�lv}���w]C}��ۡC��@H\�n�&}����3����S��g�97 ?��(nt_w 3}O�ƫ:�5�F�j��zj5{tq%���c�.����v�_䇒�I>S(ɡ���}�
~s�[8l��A�a�����w��\��h�dF�V�N"�8W����n#�����*�0���f{i�8��<����1�d^һ���2s'}���`�eddf�~֡������'|y~���[~��� ��#� �ŀ��FjNf6F£�Mư��~�&f�D~���Қ��̽R�7��Yn��p��ې9b��]���N�|�}!Y<�����o���9nA�\S�	3�r�3��ɎG��8���zS:�^+�3N<%#+�>��) �`��wF�o���B�`���I�3 bG����Y2
����\�COfC�c� �z� �U�t7�'���IG��Ar��ˏ�B�	a���&#�~ǖ� x5���Ϯ�=jbL��H[A�<��7�o�n-���������ڵXz*wQw�D�0��:�M�*�u\Y�޴5Ѷ�A��M]�S+%`u����ZNR�
��]���ъ��E�-^�i��f:AE�9�'lʛ��B�Q?�kp1y���ې����F�#G�&:��[��il���S�m�T7���1�W�~�Ҕ�
����~����*O�۳��aE��������U�L��@������]zмJgz���q7��U*8����`.��[I�w J��@6I�(��CV�^�n�H=�y�]���1o��w�z19�Qdq��3�L�f�=�^De���/���*�40:٢[�
w|G�#����C{柪��I�G����6"z�?X��)�H�]!ji��U��X��gˡ�ό�%߮�V�i����	9�9�Y+���ks�,$EH��4�{j߭�۩_�L�6�]?>��y������*
�a�7F�I�KRi���ʋ�{�rT�6���8�v��g�o١�O
1�K<�%��`	�ڽѣ��`��Y� �����@��!��<���w�(� ���{%Y��{`��^���g��Pk���R
��kS��=��ә#Y�rR,X�T�h=QQޱ8}Y�A�n�x]+�R��]1�r�bP=��V27�z%���`P��/�5���T ��Af��i�:����O�{6�ܔO��n5��c(BTC�mB� ,_��]�B�҄M�Q��?�$�5ҫ3����+&�Q~F�h6�?�v>�u�<�{bCʀ��=�M��S�HR)�����A(?�5N)�Yv�y�*���ү</�@S*�q��-M�`E�/2%'W��)yF��I��l�[c�;澥/�1�-w����&��tm�Ļc-$TQ���08u����@<S�!����2��o��'z�����8��
Aj:�|E��b�^��oxXڹ���4 ��"���s)F-Q��7�e�)����ʹtq~F���@R���Z!Ph'��J�\�,P[`�:�X����?�hg��(I�����,�jN��3` ��b�i�sOՠ�5�ƃ�21��`��D4�%���4�����X�����K�Q�9|S���3�8����g��u�'�<�+�X��F9'$�fp?�t~+�+g��S�Y��/��4�� ǂZL�D�Vggeӟl9K�Sg� t���Ӟ�׍h����E���Z���'�,�𣢣P�[=��3A���|�q�u-gц�q X����qI���_��*�8L+۽a��8��,X��B�)G��O�)¯��p���05�����}p!�LZhMd�!�T��-B)��X���a�B�~ByQ�Y�{�`����p�V�p�Y��L������j�{���h��e��;�g���8�|2�W~�`x�9-�h���~Z�yrr�<�l	l?����C�(�L{�0�UL��!�mRl� ���ou���=��jSm�d<��s�?
;�,8���7pp���5W��9�����і����)���]�y�]�K8�1�PC�A�R�e͑��*/�����A����^$�+�<��!8�[J8v�ڰ<��Ｉ�x9)�
#{m�DJ_�bv\��4��P���������Sxq���Ť���3�x�U{|���u����ʟ	�8���g=�ѝ?�y�p��A;�j�����ְ�^�9o���v��^�	������*~¤���U �J/�Ҋ�ur��P�ϸ��q��
	�T#ў\���s�e��������Aq��P�����U�k�^���<�/Tz�K�,��uVI��D{����T�/{�|?���(������d��@��r���%����%��� ��l�/f]���s�9^Νm�O���e�4v�����ƽ�tظ!�.,WޮŤp�q�L�x��o6K
�oK�B�&@s��,c!#,Ŷ��E5�|L/l�^����F�xJ��ܽ������� u$<vG�p5�#��@��@���$@B\g/�X����j��)H$����`�V��D��a��<F��9���ё��3�W�k��miwh��6{�lm���-�,ʤܤ�	���@���Q��`���F:e�2�qw^���tv��-�O�H2�2-�\�	1��̎��F��jM,y��bZPZd���e��֯2���D�����D��P���¢F�c�����ࢅ���*5iы���z@w�����)j;	�#������Ni�o�2Q@��V녬��T��P��et�J���ΒL|i�*��f�R��@*�e�P湼Ծ��������-l-�,���3k�Bm�W�cJ����$��8�"oU��\5��F#.y�,ö�:�P��c�*ʧ)Z9;���M�x���rU�Ȯ԰���VlNǝ�i^��V�����q�,/������܈#L�Lq�<�AєL��|�6����}�v�r;��J���q���\ʄ�OI<\b��f�҄CV�\��9w�V�wi�}��x��BM�L,=L�|�%��ua��<�d
]��dA�n�	��m&�O��C�Lk�s�YK>��T���½r_�f�*�Q^�7�O#�v���]%c.���5N� S<����4`�h���0������^~�w1�0��O� dx��T>qĖ�^�;/��;�IKH0���UfWx�QR!�� ��}� q*�C�lI�J�Wۼ��
� hd��m��l+.XO�U�j�]�l��~��Da��;�+�|�G3$��F��}��4��D*����OVR&���Ep�Ɣ��Ϫ3�D�����3�Dֵ�ԟ�I�TX��M��2�W>s.��A69h������[se�%���4ᩏ���m�,�����Iw��2�8���ϛT���N+W�BY=֟F4��-o���I����7�-G��(��PZ�}�W�#��}���c�z�=鑑2
�QG�� 3]j,�6�	@T�M�����`�L��$�u�I�A ���KU$\�>�1m�ء��w�!&�m�3Ag�d������>�|p/@�MfU���d�b�Ζݨ��w�/����Ͷ���GH���0�w���v	Z2$�u�;מy���i�=��1�־� �o�x�K^cЎˡ����K\�6A}[U|����%P6\>��4��k�y[I#}�V9�6T�/KB��}6�H��W��r�4�qQ�Kz
����p�h��5J̻�YO�xy[@��� �oҝ�~,��a�dU&�A�H��`���2�DN���Uf����+悻��p����X�(��u��8慈����v�h��چ��/a����խj�|�T�Pj'��u�j�ؒ�F��?��E���]H����E��!��#��F5�<m��&_e�]����w�r
��b#9Oz�0��ơ�'Č5Ҹݎ`{���y�k��[�г��dm;�D����{�zYmu�������*�/ie�5_�eٮ5�3Ԝ��Y��c�m�����e����`N��i����-싃�G��,?�>��l����X���xp���/*glH�ԑ��t�j22d�F#��a��PC�����
*g,�&<XGfz%af�mQ�o��J��Wg����^�
Tcv�@U�#of=N�b�7H�˺sׇ36�9��s 7���� f,������z�HE���H���k�]�ύ3� �w�`%si(�������N_��h��)0VЪ����&�H���`�)�i;i�$�:�j
U�f���|fx��Ao�#m��/�u�r�di���p"����XD�^b|�#�4�q<��
�s}7\ٸ��'ߊȪ� 0䖳���~��P���HO���ۘ(��*�o1� 4��+
@aK�#z7^���p�R�8?ꃬ�A���7jn'T���	ߴIjh~����ug1�������3��Ru2s�^s�4Qox��Ĥ���R�~����4pu��u���vo�'G����b!/N(6a�I$�B����#nGV?��p㜞:��ғ���_O������!k4��q:��)k�W��eU����Hz8 15�l6� ��F'��]�*�%�� O�g�����=�*t�֥m����4�r�l_����8�Zjٲ%kj�����IyPw+�_�|�TmO�rȕ{ȍ-�UM��\|sę�|)z�]{��ŋ�ą�Y���u�Necl�;��+��צ��^�_Q[���?���tt^����:�#}�XS��My�O�KG ��1+�	�B䐵b��q�$��+�S���3X�?Š=���B�Zj!�-p�:���8�H@����,ƞ��_��o��AL�ai����bHe���P꺣��
������O:1=֋��N��WF��[%�s���{џ�
3�6��i�k���^�ӓL�
�ǎX{]ş�@8��(W�HD��\������^�,+�kvw�ɞ�|�awrJ���R�?6��U*�=���k�unl�s�{,�ǄlY�L�3(��ی���!��Mn���&5wY�r� �%L��!��>����Z���t�=v�͐�@j��Ή'�j%���[��i�h�d�	���0��|�ѣm�=�s;����p5O���*aV���fb��g�!�i4�	�""�1�+�<�����w��\��E�'~u�,���4=F����,�������Y��!�As��cyE��9��"[8Qd/d:{[�P�sq�:���]Z� ���u��D�;����:����iǁ�31��E��~�<��nɜ�v�,'6����OL�t�'��Tq�Do|@0��9klALnk�6�:FJx����Nヮ�Ɔ����Y]>�f(�b���:�D�d����g�����G���9`��#h�Pc(#j��t�"����[�����0��-r`��ݩ��m0F�!��a���p�o�t5��Gu�k{���9��Y�Y��4҃���GR\�����J���7��h�;nA7�(�`ͤ�l�L�u�
�O�F�m��/��:�z�c���qw�u*:#��e��s�0(�/,p���m��_����i�%5,1��ܤ�Q���jm]yE�!� �w��tw|� ��j��#`Q�v/�|�W�\*��9��@N�z�U�}�O�=ݒ_���*��<C�?2�*�]��*�W�����G��L%v��[���z�\|D��E}��dZ���-�������&��ǟҪZf3vp=^� �~o:�`��=��������Ui��m���/���c�_��/U�(���d����V�Q��젠�����w���'Ά���]���]�la?H�	��u�BAQ,w��Dx������N��<h�X��f�W��3�������9���*)>G�M��?1�y��&����^��� QZħd�o
�0���5x��}9�LXV��<�7	W��_�(��G"<�*� -�Mi�v����~�X'"w�/mkp3KUֻ�qyO�qv��W@��"0�&F�N.�$��;�g"��7?�Xq�h���,�}�IC()��XⰧy�����'��)��J:f	�d"�
����n�~G*o� ���Z�"o,F����7�5�$�2d�1�<��(�D��t�y��\�%��1�-�~	���px���?D�1T:p�l�s_��v?�	�,��j�䣋��.�c��%7Əb��1B�z���7������f��\��f��O��������!�~�Z=��iH���zhs���Xx�3�a�Aw���E8��M�O���
���#��ʎ�}�-}�D+�+ܷZ�s/ �#���L�޹��Wşq�:a��-i9�E�*FA�Ɯ���._�������DN˭�S���
�u�+�v�����Q��k.�rJ�2��Q�K����9�����\]]f�&��%�!��E�TI\�B�H�%=�&>��z�:�?�`����xmɿKze��{��$V>
��dõ��m�{=0������"�+�>�c�a�g�m
��a��іn	��,�O�����!d#��7m��'�-:B�9|�:͇�|����N�UqB0��dȎ�c�)XuXlxVHYEB     24a      e0Ms�秛s����
3~LB��P)��� l��5�	gu������>T6�2%��*�ӆ��Fm+�>��@9�<a4�Nt����#���N��h�ݔ���t�8�"L���%��>�8.N&}Ђ��*k�	$A�s�-�k%	DZ��o���?_�H�U��`&�j>�zZ>�ӤE`�ƞ�K�B�`��C����9,16^x�^:�]JD?�]y.+�1ݔ�R����W7�~