XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������eb���:��@x������ 愼����1G���uF�s�K���5�G�Jz�W��m
�b�����$ V�v���0찷�6�0=�)���e��7s"r��L��k�k�J��V�n�I�_���e����z��|Y:I޻A��@�$���0�|*��e?�9Ԟ�#�敄*�*)�j�_:C€������|����n��s��O
8B�Mp����}�!\	��*�u�n�����E:B#����N˫w �)��Y&N�N�x�n�p2+©�C�n�q����b���?�=�)��e�S���>��7�x�̲Rhr�����5�b�qv>�_!�Ӑ� `���>����L5?��p�� ���v��Qv�L 'yfd��f���h݃Z� 7o6�L�W�Í!%�o�V��_t)��ى��2L!:eU��~����c�",�Aa!�`B]_8	�i��w���U.���'�ouX�%�9�5-DYq������@�;��T�?y1��(Us�k�Q���@0`�q�:�|B%w�� 0f�.�g��Pb�3 ����N����eo�A��{�{���~�Za/�)(�TF�5�K$�â��g!�d�:�g ��%�Ƴ���٤����A�����[K����Yt��i%�CW5%*4K�-|�4�X�a�e��,�/��zo7eI�����:h}*����R��ڃ����
�y�*�K��|�{�S�����p���O'��En���.j�u���/���XlxVHYEB    157e     760h����k�t���&�?Z�����3�L)��1:
K*"fq�§V6�2	(Þ����2x�Cz�D�ΐ>	X�1�?T�R��,��E>=s��'M�΂>S=F��,��z��y�T�wX����ެ^!��ć��-�-E9���LtM�J��o�>!Q�H� <�� @>��xw�p��Cf��������^8��ؑ�GȎ����#����G� ��{ϡ�c����;p���͊������D:�X2�2�3v�����/D�Jb�$�}��C�n����H�4�G�}�w�!��{�ă�i�q���j}t�rޛ�Iz�,~���;b6�@~4�����B�G	�]/�7����L[V�X-ܣt����k�8փ�%��M�v1�㑩�)�~C��y��|k��S&�ɪ�d`)�I-x�6k×}�2tL����j=Tx�9h�B������#����;y�y!��ch��f�\ �X�A���d�Z�AG'�����m�Wq��zs�64���e��:U��h%訣D���K��hjYs>J"�9�#�����(z�m4C�ƲT9�2�{]��6	 :U2d1�w�a��7Fj>�B�����@m��G؎�k]2v@�"&� ڗoO]k��p>]���1r�\�u�s]���/��"��NX93�(|4�}��=G8ޔ��c\�޼���̏�Z������">ڃ�UN��TO(�����B��� �H=�L�����Ӎ)/
b������U�p�4����i[/��{ΰ��qm�B|�p�$�r���G-囙5��>eь���]T&B�}��|� �Sqx��!F�o�rӳTy���v�j��̋`�G��nY�x������x7p²��Z�t` t_͵8>Zv���YZ�m�:Y�,��^�q��[3��:��ĘR���s�:M�����=�N5VۇQ�Ovسl7������S��
 ��w	]�ӓ��dW,^��]��c+ʼ��'k�C�|Ly1UB�Kl��m�����cH�X-.d��f�UYׄн̈Ig�C�_1�{�L��Ab���WKBk	�/a$j>V�M���9�*��&��H�`����8����	گY��W��=p:�#��vx���X�ł'�ig�I �<�ܘ. �WR)s�+2�qov�=�S��ZӀ��
�3'�����*گ�Ľ �R$�K{����~�Ǯ�ÇPh�+�%����P��5ҹ5#���ǖb�2�[N"�;,2���O�3���h��B��1s���M���s!s�u�Dq�
NG���ȥ�?k�/hQC�3���Y���8}jԪ��%� h��^씅L����h�h�@]Z���x˼I�m����{�G�g�S� ���g�4X��GQ�a��Ʌ����0�T��pb���]������v��{�=�ͦ���}���,UI!a��b�HE��`E�I�N��l{R�z"�����`l�K��1�K�`r��<�����h�G�5��p��,ް��A�u`��)�يb���;!�|��]�2�q˥Nl4����|^��O������H����F#��V�H�BO�Ak�;�ćUو(�nGl�#�>i����"*�+�����\�N��GW�d[��'�[0�h7qk�@N>���~�`+���@�1k�W���l��-|oҪp�Oywt�+J�@��G��JG��4-��c��,򓵷΁���%((�&����YTֵ���:R�(�=�3#5A99���Ρ␴m�`�,�0d�1����CZ>�@��BFU�K#��4�v᝝Q�~���eZqw�Cp�� ����-�RF�E��U���I�=y݂}��`wT<D>r"
� �O��i1��v�>PF��X��^e�