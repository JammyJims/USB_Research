XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7HׇW��M1��w���"�K=H��m+��@{�׿R�*�=�p��߆��_�m�禉ۣ��iky��
a�K�A��f��e0���lo�~�p�֐��p>�9�s� �s9�mM�|��!T�B����L���!�����Xmū��;�(c|�&�-�fs�b���o��O0�+V�c�seQN��r��Ԃ���YGT����rc�
R 	�TF���Μ@0ڡ�v��Y����	6�i�tc�����x_�����7sd�%zv���w�,^G�¸}q�q�;�I�dʜGe�G�k�F��%��U��xn�P����3�t�]� ^J�ѡN�!Pl�i��ڪ��(�D��qY��/�6�~\DOi|kؔ֡?�L~����D� ���-��ym
�2%�%�rt�IL��Q�(I��������򳄨�	r�,g�\5��"�+�*mm�� �&A��,oH��G53x}����R���d?4u+��{�me���H��q�K�ᘽ6_�3u����C�Q����Y��c�����+Ɋ��1��n+���Ly���:�����|����˼�і� @��%8C���r����X&JS�s߀m�x��ϟ,-H1ʻ�h�7qZ�U�a�<�~=	Z����h,f��g抒ARh��O�B^l�b�ډ�������F2��MTr����:	��5��/�;ܵ;'jir���)��B�p��W���F4������A�%�@�Ү{�b�1��J��;�}S�RXlxVHYEB    fa00    1730�|�5���|�?�X����:�M�e�f2LRʓ�A�N~���U񿠦��rH�Q���P�������v��F7��D/b�*?�7��r�'��'��osӉ{	<B�x��[�`�����O��5�e�5#�}���G
�����$�D�H~ul[ܜ;U���5�8�^�5���!e0�w�9�a��Ӡ���B[#��u���E�&�����sܰf���A��Z���8��q�،���h�q�=�q^e�������"�]�����B�E�7!4a���EM]#�P3-��L���ƭ�1�ʶ��[�>wX�� �ĪP �����[lt(۹�J>�!��%t�٬�_�'r��c�`�/h�\�VȜJ���P���K�3Ӳk/�fy+�b�K4���?@ɮ��-c8y���ZEc)$%��	�H]h�G���[�lA谌�N
�	8w
a����M�q��� Zo�=��Q�?��0��^�ò/�&8��,	{G�g��uRq���o��q���\^���
�T��V�-lkc�+ȫ��;	��:!�Z��*�d0��5�4y�M�1�,�k�ʓ,u ����w�Ҽ�cvz�i�E�#��K�b���[�6���3�S�5Ł�9�ϯEYC"ϾK1���f:U�Z�	�6zF=�O�2.P$�k?K�rPs
)���$k�9u6�tCD�Ξ~᧺��dQ�Ȱ2��u7��A�ÖOf}ӂÇ0�[�آ�a���cD�}���)�uDt^���ؽBW�rp��#��d�	�/�
�<�[<�E)K������)c��<�jp����~�B�'�B�M
��k�����WH���6�X�eH'����^?�p��Iu�D�<�����3�_��"�)V�A]yf���͏3�R]���uL�j�G�b�)�1%��V�� ���^��"G1�=�rv�2���k��f��W�#�U�Y��	���cCϛ@^�"�4u�,��]�A\�sٓ@�'ؕ�O{�r�%]	3���H<�O����򲌱��ʏ�s��Ӛ�M�3m���W_QX�c��COkB2�h+e�ㇸ�ۣ���$�s~l�C�ENz��3�l��X��,���������M��k�=�.����N���70.\O�}�Y'Bh~}�#�s��}d�j�@����z&�*(�@'
�r# ����d�T���8?��	o||� �����9S�0���=O��F���-2f]o8o���]��o��y+�<o@�V�y�2^/ʺ&�Xm��nβ�ݗ��IY!�n'��ŷslX:8��y_�� ���8L�(��������޻f||kOOO)������5M�Z��]@�y��-{�� c:�,k�Ðm�+v�F�3�ߪ���;��W��2��[�� S�*'ٵ�z�Bane	��*��y���3*��'ja�2�dHa�쓦~����(�F�+7�Ze�\����.L��e�yo�P03���9�	�h�z��r������gO�.W�GuiЯ�c����H<�1��DiY�r��\��זJ�t?w[�ĠM�n�fg>x���'��FJN��xTD�P�|��=�lf���� �=����9�0N�w}��%��!�6��A��Q+�Y�ӓL�K�Qe^�ZM8?$��D}�Zw�%�E���BHS�k"�Op4a_*�g��T���B�rA�"��	!��Ⱦ�*V.c�^��&a��>���-�~��͝�G��G>�Hx�7�J�5U�S�z���¦J!�V0Y%�wq �q��6���;F���s]ηY�:[Q]�&�F]4���M�F3�WQ�W��~����,�r?,�m�E��k����YK�$WeA@�{t�f��|��#@Oΰe�����^"��e���c\�9�X�<H�ȁ�(��2��R#c�uI�s
x�Xj�|��dI�D/Z���.I��q�G��>@_�����`�!�^�أ,O�1:3�� �z�d�d����j�����HۢTE�l
�X϶Bv��jf"��0��3J�% +�d�	���ל�qV4
��^���K�[�����\?���q�b4��L��'��"�`��:�6x@]����+���w�L�T����`x������ʜM�ӳG9�om]nܧc[�I���s��Y�o[��:~�!�������}P�'�����51�!��P��	����J/]A҉(�5G5��F����uY6_�owb*\/�Q@�ȃҽNqԴ�$�SK�}������d�p&��&H�7���g��-Hl�xæyL�<�C���ޖ��-@r�C���/ݖXbX��;�Ó&5���s��&�r����},Sq=P�+���kѱ��i�$[�Q���,$�k�ɵ��	!��}l���5A�Y�[V{��Ɔ����y��pl7�U���fiI�Ό<�P����C�^p?����iR9s��$^�����-��ؤ�,x|�GI��
+E�3g�c�6;�5Mtՙ�p j½���e�J��dϰ��R�a<�M5��P<֕�+�x0����"��87��ݚ�����s]x36â-�LE5�P0���#�w���u���	�r��D�nl��x1W�ɘ��1���^�b��4)���3�
��x��֤��H���@#:ot�+���sg�U����B��vS��HpwJX+p�BR�C��JtF3v�P�O��O'��^�q�c�؝c�\������'<�*c8Vk]��D'��Y8V
ܒߓ���.�~%H={rK6Y�^��&�1 ��3au8jV#��'o���K���w��^��n���Yhϩw�a�umB�]�����P����H��d�&�X$ޕ�h��6��8��:�����Uᔷ��%Z	����B;�>Rψ�%%��q:�Ȓ�Ҁ!0��`���_WǬ�5e�~+���Q?��i��/��<̃((�=��j�k06����s�&�b�?2ೞׁ�(��
�o\\�Ž�n�`�;'l��rY�L�e�v����|�ڟ�\WU�� �Ow�;y�oo��nhi:��QW���C���́��RD�B��͆��w�.�(W�<�%�$#o�lVzM������m�eC�=�ҋ�'�oʄ��r�^�kvHQv���*����`����?�ɴZ D���N��(kf��I��޷�X�N+|��}�|���2�4c��9������e�QT_]�0�c��/Ů�˓�ͨj�2��|r��l:�g��F^p���d�e�d �ǹA�:3V86��W?4����m5�{�ە��������e����;(�@�l����n�Len\���e����5q�ш��./��G�
١{��4.���0�{r{�	z�)�.��􋇬5�!���}��K�B�Bmj�Ňl�]��� D�%�7D��	��ד�����6�� ��9����g��M�KG�t&�jS�jV�s�}��H�T�?9�)�a�"���6[������L�+�1}������
����*�	2/��`X�����e�ba�dGW��cr�8ʚ�3�6�!2F*�˧�Ó�߀w�L��5$�ۿG�FуAw l!!�Վhy��4���w'����l	��i�U!1,�<�(P<��!��zBBe�ڈQ�,pw�b틚���Pe�P_t&�Rs �
DmuQ�ޔ�q����I�LO������PU����[�SK���SP�%$��#�\��/��|����㥄�)�Ϥ��f��~���x@��H�	������g�OQ���&��Ҝg�)"���ٱ���ԍ?^[�S�hO-������yh/�F��K�\��@�0-'����	���Ft�>C�,q�3�6��,~�b����a�#��%tm��-w�j|"I#��.�C� cF`D��X�PDﱁQf�9�H�B����|s_΢����X~��Y.��ڸ5���+�MX���YurbJ��c).�� L<n�p��R��#���/y���	�f	ѝ�t��Ҥ��K��pF��3=����\��y4,7 ��q_�}�ދ�DRV���&��ѽ6�-���n߉�����mmu��E�x��*s��7қ�&a|��� s�S�y�3�։2G[��9��~��~�=�fK���9Nw�F`\_��6� E�g��-d�f"���{���[�U��7�2�]vf��8����8�#
�~ĜhXͯ�@�,��s/���<�G^C�*_�.=�`���:z��ռW��a�CW�ٌ�*�Kc�4���$8�-��@^Ӊ� i̲۪��k�k~���e��qw����u�<��P��M`�$q���ɤ9W�������]������x���=Tަw4�-���M�X�r�یe��=�!^��?�^B��LnE���
� lq����x��η��f�
�L��(�e���7o�SoG�Ce�-D���b$Vqw��DkO֮��T>�!L�D�8�B�0�!�2�U�A)���²>c�g�O^��*��>Z�!`���)�����U���51��Uj���X�ܡ;f��:��$e�3�-�b{�V��[�	�8g�\��"���Q���7��F��� �?_dl��A��;�YoF�}bӓ��@��S��5��KfYo�n�7�cs~p��*t-���C��M?��T��|1�8u�;�V��b/&�#���$��cw�<s�[o_ڒ��V����;S��q	W�cX�H4r����Mgލ��҂ѱ�u(j��#7�k.x��4F	���������׮�������� �ÿR�!��t7G\+�*����}f�C��v���I�B�	��!=x�*�!iD(a�+s0ë�*�}���HT=�T����X����~��W�P�(���,|E��<�«vu���%55���� ���D���*f�Ǥ�6��i�&�J=ej�+�-"�E��i �Ҿ�CՌ:���P��܀#��Ϯ���3Ҟ���+���$~A��3,O�J	��j��<�*�o�+�h����.�r��}��hh����M��J��[<{��S��6�9�7�qؿI�rRc�N��&�+�^|�I>��ٍ�,g�f�WOU.>.R9EF��	-��^��$��?�*^���ˍPO"��C�a&q��W��g$/8���D7�@������u՟χ�1�Ens+۝(/0X����]L�CwJ�2�|Y-yt2�>'hbY�^[]�k�-&�I 1}�A��y��]��t��0����,ͻ.u7U��H�l����1�
�=\ ޝ�>GPM�J�a��-6ԩ_!���/d^"�̭ ��@�s��R�=R�he���y�=�Q����fT�u��Vn	bj���#�U^�p
��_P#�~^ۇ��PY��I�K�S��ew�O����,o	ZYxQ�F�5�n�.�ش�0�ʚ��?"��h�h�ML�aB����d\���N��� n���sw#�h)�"��q�W�Syş�6�ik��#������r�����2��װv}��#���VT@^�'!=D��SZTx��D���
��Iv3~���>��ҳC&���P�)�X����=&�Re�����0*W)��CU�B�O��}_l��䎮�Q�,ԋh�[L����aʣ~B�ˀ��^�FM�0�ĥ��8-'�����`�g��	����f��:�ү��5�EF���i/|���C�������E-#���Y�i~ӑޙ��JЛ-A�Xp���j�2�}�o��޹��-[)�����pM�U>���cۨ����wA>{��#@dPDu蜻h#u�U��9��
K �&)��=C�@�B�d5|��#F4ޥaï�k̼��wBlXlxVHYEB    fa00    1d70��<���#v���g:s��i���_��Pf:->����5 ߵ��4܂��&c�� �do�����ŞST	@����m'���C�OE��M3�|�5���ۚ1�����F[�)�T��d*�zc��׍mO�6L;ua�c����l�R����7l)�'��~�[{��&�,G��Fr��'A7پU�DyF8��V0;�F��`�[Ecm��N����;�������V=�t yI�]��uH�!? 1���"t�UB��ЄQ�t0���u}��;�7�G�`�|���*�W�2ե�v۸f"C�����=��y��z ��H��vxÍ�O#E`�"�m׍]�����%���Y����>�F�qּ�P� �`������܌���Ϊu��l�δ�M�j�$�S�gaC�Y���^1X�ږ����cub
>���I��LD�1=�El��1:u:��1�����$� ��x�h�5��$�6�@�`��n�m�`�g`.��E���p���X����P&�g7���y�m pIG�~&�
[���x�Z-`��'�km���Yw�b�Q�W��/���=B�>$;�s�;� @�����6$��g��魈C���}��vݵ�s���[:`�0��NAǇ���xFiXA�'x�>;|_T1d�9���q�v�`�{w"�0�� ���'5�ɒ ��i����"�c:������)0F�×b�(�l�'W������>@����8[F7�PR���3�$��pdu0G��������77U��2�'�K66�?�)[d��b�03�����}!�q~(l��f�q�P��ԍ.Ż@YX�����w�5���8�3;c_㩽�8�Ӣ]�zU����T䱤���g a}5���F�_ ��2�%ׄ?-�9%'�߅?u{��7�T�I�qԶ�gUS���h�Mu�ZY���/��Ⱥ	�H����L��K"���O������^_ea�vJGе��ڸ�>1W�&���v�	�`GHġ"��+K^OG��Kh2U��(�> ������&ʅ+<ER �!���]�B��������|� ��w������;�D�>��T����@nkʋڇ����wT�`.��7�!;��a/�}����l���,Tk�鷮�U���A���g�Hr0��?����陜�RA]�$�T�~�[^Q��B�a!8�$�-{�bN�Ge��'�Y�W+��*W����I�	�+ z���oK��x�@�u9В��_r�����Sl��w��n�_ĠQ`�-u!�@϶�fX��UPP��[o�蕚Ġ�-&�W�cD��@��ɧ��Y�I�؂��a2���VZ�'YU��Y:���W���ɑ��)��bzSޟ�<���lIIq�}�xs[|��zL7��i_Oծw���s����,:<��N� �}�%o?FN0����w�r�a��#������4�(Umi��	>�i6�`i8-�!̲qS$�������r�2Y;Qe?[ ���S|)�^h���M��Qy��|�Q��vJܖږH�cR[�4����0U>��Q~	ְHe�ζ*���sc��3FOP����%1/g�h�΄KftU�x�_'T�¨����z÷����������ƃ���ҧO�\�vk)�[8�կmG��!�D�^�³�s�3�0��uy�� �+�=�J�[�:��Cm�c��Aƺ�^4�Y]�8N|�8���K�î{J=�<!��Q��Q�IA����?�D��)hxpf�j%YJ	�h�!ѫQ�����7���b3
q�@��H�\;�h���W<R�u<�K<�f���āH�����Wv�_���>�^V
�桔Ÿ�*��r�ڃ�+�����i�WǿS��Wk�M�6�1f��nW�f�bi'EDl�7��G�-"j��R]�/�*;ܸ��" N8b�X��"<��	.�o~�� �2� 
ܢ�w2^Ә	��άq��2!���(�JFY�� �!�剂�D���ǸZ�`��p/��b`|��T���Q	zc�l��ta�B�2�!;.^#� �B�1�^4�wE�_���'}�n'�B���A#KO�����f�o#Vj��֣�#�~~�R���rS�2�6v�?�����_�!���" ��{�9�y!b�x ���b���n�/�X�쬷���>��j���DW�<i� m<�'�W���IT���v>qQ*�8�X�El�AȖ�a��+$�C�Ѫ�뮊���(i���J�0J��S�a
�}[G�:s�����ԶY��bɁ��Q��$ʸ%^�QgR%�4�s7]�Fk	s�ۖ���9�MϾa�wuh)�1�ղe�8Ϟ��X���>	�3O����6�3ÿ��v����`�@��W����y�/SGfY�}�9�ܠM��b����M��p�,L��� �_���<e�[�/�g���T;C�lP�Ŝ�(Op?w[O�N23vk.&<�Ye,���	d�y\0K�ÁC�I��q���ݥ�����U��䱜|e*�J-�`��n܁�_(9	B�|��B�ͅ/���6�\���É~�?]��.|V�>�_����B��׆D��q�L��x6��4<O%V�:��B����G�$&_���,Qz�HSi6���l���Tԗɠ�3(���VRå���~f��ńzW6���.��k�'��z��N�R����b��;��rS���n������6�@"M�ι(g�yR���0>'Y��'�Ln�k�~y�'1��W��q!��;Hx⺧-O�����~Od�NF�iI��0|I��y�siۊ
�w�-��2���CgI���}hZu��s���<.�SGe�`jv�&�^���ɕ��Y�=��F��µ��Wh�������^�M����<�bJ�S�
���|WL<�!.��%��!�7r�2+�'Ʊ��S����U���}m�a��!U�Ǌͽb9�B�q ���p��z��P	��+���H���{~�����F��`�?�:v�J��.��������ت�[ME�T�2�4�X�|��U��$^�m��pG<�&���V�nH�I�?ֹ�7i�rZ���s���k���;�`��w�w-5��&��9�i/V'��j��%.��4`k���?qw��hAK��G5Y6��y}b2ը��B��_�8�$���L���J���������eJU���!�.6-��,0�2�-R��k�����F3[(�G�S��ɭ<z�ҳ�����E_���*����e	.�!V� _�s�3�0"��x?ۡL��9�<L���>���i8O
��\]�c�[��&� m�X�a��9Q��'E�47��5���h�2S��D\`�K��0�M*��۰.����D����]Zx����~�X�#d�U���QZ�t���������)Ep�(�����75i\�\z�o���q��ꬸ�J*���u���/[�t��sw�aۮ�|>�q�¨��"���r��@�E>�QuB��yS���B�~'��}�	�M������2'��L�t֐X
�ܦ�S��3�iE�vd��%�;���ão�#�Hem1���|C��\��eC.\��m��1*z��[/����R�|���]�g�:ɏ=	�2:�+�Y<�	�v�J$�����!1INt������df#iVy��
��y�M�S���o�{���%PK�ٜ�Y�v`
h&�x֕��,��G��V��S}��+��$L��k���F>���VF��F�k�_��%���ٗ�� ����7�s^\�o�d�� ;���Ɋa���|�):~b\��y�^!�'5�CZϧ�4�&��̃���<ߦd����5�����3��i��=G�`�>t� �/��\d�~��-� /���+�H�R���iM0woo��@|����zdCgȨG1ь�J ����=b|��} ��#d[Κ5�s��e�#����p�X\�[��%A�mFs ���E6���_�cR%h��# ������s6�&���R����g56��R�c�<~��o@b��[A�,Ն��_���	+H����z��c%q�n��G�4��zct��h���w�g�0�X�`��g�Jo���f��HW�k�u�"�6��hj鶯V4p����}˦��U�n��6t�r�fͤo����hTfwq���,�27�-���(�I�POբ2�ʋ 2��A�QEK(�)P4��&v��Qv�#�H�ț�YD�׌ڢ5��Ɵa���q��i����.��J�}(q��{뵭��PO�R:��V�Va��u"=xu��D��?��F��5i1��S� b��-��ߟ���"�|I�G�'^�P`�A�/��Z�&���6,���4ߺQ�3ZXi9Դ�հa� a�7%��S���>h�Y��Ro=5F�aQR�����}"�X��Q�]�=�� 6��X��	���	����Bk۬�e������g��t2�F1���l2f6����@I����{��^s-� ���ڳ�#�|\���mm�)�\#��OU��	���>�v������3�}��l�cz�|5G$h\����:�&����@�哾�U�s�=G2�("��>T�w��m�I�N����lf���~݋�?G=��RlQ̱����-���-XK��-	%�#pp�ջ��gl��)M�Nq&�Mw���;i9+"�@[2P�6'e���:J��c�b�̌�ϫ4&� `����C�?i�-����1c����ȶ�L?',`uidk��̭Ť@%�b��M����%y+��B��]�+��k�(�_XQ���Ҥo3u�^�Ӹ��L�2����Ѷ�N�V���L5N�ȝ�-��YrهU:yA��,��
t�~�9�B8%s��s��,q)�"@h�Y{���f{+
U�xP�{]W���l�c�`�+٥��e�	>*{X�s���Oh���X����<��_�U�X����MǢ�^�X�|e>��c�F�����)�-���: ��+T|<ǝ.����d��NT(��M��/o���>��C�*TE��0a�&'��2��]�Vg"�P��5���c3�; �y��ɝ��h"!��c��d9�|�Ks�K�љ�d�)3����43��~X�����ؼ�j�N���<n}�{.}n]�mJ�q�;�4��x~�Au�랈Ӫ-������>���*���Lvk�����;�7��RY���_�O19+��l�0�u��
s���	���ζ<�e>�a�6r����\U��{����U�������(/˦����֣�'nz:�Q,����M0�}�~�QQǻ6FxH'��׷��S�HT��|�=N1���z{F����$���_�l�g�Q�2��z�]�]��{&,�r酼�NL�v.�	Հn��Yu��K|s���&�x�z� ��n�9� y��ќ�fj:_'Y���R0�9k��a�#��mҢ�I����\5-I~��wfP�w"��*�r�J:�Wt��v��.�I�E�H.��J\�ʃP�����fn-l�6L?�m����>*�d;#\l��@Gy�ƽ��2�y�J�a6��Gzc��m�Q�9I�8�����0��7�'���XD��~ ��� !����f�6��C[�ϕi�`��j��(��:*O��x����$�2�E.��)�)���s:$����.VV�\?Xl�}�;ܪ��7�:�~��}�x��>�����p�I�(~����NW�D9I0+�ㅟ��3�L��|�[bӿ��G���� �Kuy=sX�����u�u�.� `���9&=k���˃��M��cI�E�"��s�ZkG�H�D86
t����:��tQ"����?�"���r�$�˷�%��:<~��i��GUx�.��s��L����"LW�7<o��{=T��r���$Dl�GPU�!'ZʒG�n�a����8V�?��4-�W�a490�~�rȧ�{���H�͠���gl\������v�j��x8^�y#h@duJK���G�L���}�mX�#���)�ؕ!j3�~�a�{H�B�A}�A2}=��E������:�	��؋)?V{F�P<��X~�Vx���V0O{���
����>4TT'�*��}�:.��n�9J�i,��K��HU�ܥ������/�A	m�~E��A�PG�H������Q�5L�����Hbm�����U�$1�"�GY D��@��o�r̄��w(���a#�G�{�}*�[ K_k��c�ӳ���m"�?]��.�⚋=�e�א�4�Ӗ���<��L��%0,��u[�S+N˕~�1�������Dp@(����>~4��τZ�O�?ݎ���O�8`�R'�͞����l 3��
N�(���HX6JD�76n����H��6��o�b�Zۼ�Ds���*�V���)��I�N�/K%�:�/JCe��:�x*xaղ�Y��˚oOp��է��/늂���UYN$�u�mk�[Y��� �@>-g�u�l��)�L���xك4LW9��!��vf�i��!)��%x@ه��c�w˷�UĈ��-tEw9�g�O�d�U#���5��pd����k��RhD[����*�x�`�2�BW�j��<)����o=~zTu������MCr��ђF�d�y� ��1)��2�F��=�"6�hl�97y6мR:�:�|-�ˉS�m�ui9:��%��o?�V�]��{�9�^]ql ���to�$gS�i��	+]TI&w��уN0��$�|^�Lku�9j�c2o.��k�y���Zm�%E�����:#�}� &z!'I�Oa�(��V;���,��!���e)�>��t[Or�|	zJ:�N�4Q&Ey�Ƹ��E��I{>��	����z##�o��/���!S3�"�~-�m��g �5�T�b,T��Z5m�[���kyB��фy?�I�z#,T��n/� ��C������*��P����^�h���z�<F�fx���Q�w�J֙h����<���Bfz����Z���]t+��;)
$�Z�����	VD��\�UkR�t��A�8[i|��J0nD�FA_<	V�����ߙ�6�b^$T�#��B?��.�| )f�\7�%5�*B(�S���Y�մC����JG6A=��"�_�cl����G����_ ����*�n�O�����t�y�@�+OA嵃9�&1�(� ��K�>��P�h��7����t�6���dQZ�i����ؔϳ�[���*`���80E�^ى���=E�_Ԏ�_C%]{�F�TV�`P �����:���'��p�I�D�:��Y�g�\�
����
z�kr4J�ã��O��ѱP�����fm�|̓B��;xN���f�3]��yT�4�4��
dA�NS�"XlxVHYEB    719b    11f0���c�ݪK��hйؽ��0YߺO����ot��m��/� ��rQJ��v�B�&�Q�	��.���HSfzP�Z ��k<C�u%H
���x�˗�1 )hve�:9_
_t��oW�0p�ۊ ����n��Jp��!�ȸ���Guc��0a�C�J�d�ήҴ�I�ͽ��l�iD���P�n�x}�(�Z0�$4�t>lg>5y�Fr� �d-��i������ىu�An�F":�(��8��!�8��P�KƁ���(����;��K��)<���HWj�����K�cf*�&�ЃOe>gz#󤄼��/�n�d�&X�}27�Z�؎�]3)�qh8
p�B�¹z�Ѫ��<�Pd�� �YF���"�,`���>�͞/����u�T;(U�M��b�Z��o�6���mk���~��:���Yb��{dT���5���>�~�G�S��mj7,a삳���w��󬼯(��ͼǐD��!�=�Y�7f}�|���b�gsJ�t���.x�� ��!NL�ውc]��z�:n��mՍ���*%]^�x[�m֞����݌�=1>�ʰH��֘˿(	Q�E3����``���H�4��]�l9����U�`��&쳠u_\j~kF�+�fq
�m�,��,���n���cS]��Z�g\Op�^�1��{s{��/C	*�N~����~s�jG����P�Z��9*/�&5�A:w��m���A��q����?F`w=���I�6^�Ƨ�Ӆ 堛��{���3Þ"��h�%`� ��@�Nl��mE�ޚƱ"��i���Y�.)���M����}5ʋ5�b��̽�E�m��%���,Ħ-b�����&�� �j���A�c��Z�Sc��g*�N��i%I�\�:����m�FA�-��u�A>`�n���9��˔���p
�d�?��՞r����IZ0܉�Ӥ�@��2,!{�yc�����8p
�������@&���cLbDN���*�	`X�����9��Rlvv��܉������������ѣJt�1�P����3��VГ����z���򙤺@�����L�3fx>�)E�����..C�����!��<��
$��iٽ'M�����<!,��ύ�H�6��\����x�Q>�.� 5��v����m�4væ���U��K���s�M@a?0�qĂ�>�~�VWĨX�R�}&��Z>���L���VÔ��E-	�Hd��WGWMa�<��<�x>R/�N����>Ua��B0��A	8
�No���YGkrC�����A�h�[=�$LW�SҊ��L)^��$��[�͛i�%�\�Kj�LK#�.ƻ>��+��,	r��K0X:2����H23�+��ѻā#�ڻ��x/�5i�"m���gx�t����_H��<M#�5�F�G|�P��p��O�aG��%��mv�u��gɗEMe��F����h��� ���������pK�؛2�R|�iҌ�eqK�k��U���;�]�m��
�[�:CtkY���{5ύ;_�Qs ;TT����ȬH��	��`�֞Et��.��]|G�8���ベ_p�ǂ���.�Q�fO�`o��9򆎩W�	���r�x�[T�-e1��>P^Q��� ��5�����"�������%���D�,�y�;�哭�4��	׋ֽ�&H�m?/xˀt��}J'������KS����/�RV�=&���0�%����m�e� ���� Ԡ+ �-V�9��:+G.+t{c]5e��Y�x�2�I_�M�s�v����IǊ�Ŧ��D�X�5�$K��j����<���]�0*��{s��3�o��a�sc�4��"Z{��w�]�=N7��BۢtoYi}_���:���Ɯ�wi\����rk�.)&�ѹ���5�1�i���	eM�&CT���7��,���wV��rǮS�p����O	�m��5�����n��Fi3�������)�/�9gO�y�,���ٜ,_kRKoV(��zWZX;p�f(RϰI�1;��r��ywe��.���UY홍�
�V�pX����ש�z�Ț^hNG�94�"=�%�1}���o��jPI�d�`ؓ�m���8|3T��+P[�̇tR(����l���N{�9з�g�{� �����S�x�=�3���F���Wh�:)~�VG�w@L$���\�e�F���kH3hy:��j�%�!�~�w���hb���u�,K���+����N2^��Μ���L�VLD��l���3B�V־Tc@���yRF��NB�L#6dO4I�Ӌ���{�pV�����VUÎ��p1����yjb�p��.3K��5s�ꕧ��7�>
U�����rm��!g�[���}�Z2�.k2N�Ӑ6��]��`�F/uPv��1S��]<�u����+yYV��"ɩ�+'P�p$��*�²��=� ���7�6�V����E�c�'0�a B�!\h����*�BO	�q���`"�x�`�N��QFQĠ��`��J�1מ�%�إ������@4Ù�%�l����^I�M�Ǽ�jؿBX|���el�����9���03y�ݚ6�����h�53��^FӪaf:�����v�W��n��Ҝ�=j/�BL��:W��A�_�|��</��	��r"+ ]��*��+�/>�ĝ�-�f]�f���U�W=?�x>�x��U1�|N�� ��:��ZY���<�N.��Y��6��	5́�Xk�u�!$;t�(�;G;�=�e.���|��!ˎ��Lo�;�+I��6�Jj���U���^#��?)̗����-��� ��"��i>�d�0"i��n侱Q<�v���]�N�tT��������{2��d��#`\E�Pd�"kh��xx�c�93�qҍ�7�W��g��A	S�2�pU����7���>}?r
;��(�^���M��M?u���jhY n�z1�|b$	"�ŻHn7#���i�D��/��iSv�8H�C�Y-�y[�n[�\��"4�g�<S�,q�^��|��̅�#1�j]4?&_Hi�ui��h�\l�jƈ샯�ʶ_�:Z��DH��+YHg�>!h$7��Q�ኳ��b���@n
Ec�(d@?=|��>���A�هv+ly�Ͷ��Չ��ӿ)G1�D�L�K�s��^�������;�Q��z�o�������o?ݙӑ
Sth�X$��ly4v���xÊ���dW9 �����wU�9<?ZE�#��ZƔ\:�-s_�^$3�zT��������Z�3��$BA���[@�����M�ч��5����?��tw=P����HH9�~8cef�K'�HCQɉU�1�d��{���0��t��&������bA��@_�|{�B!�o"b`���!F@�s��/(t4�eExs�9I����Fh��%k `�%Z'��B'�(���c�Lyf�7�nGWF���%�h|�h�T%����N·eb0�GMfҰ"h�v���+�%��ԍ��I�_	_�̆0�etL(�|�~K�4�RO
��?]|����:^{�f1��ȜM����惓]�޴�M��O2E�L��yr���,oGj!�DQ�>�9����,��7Spfm�tWX&!-|��$~|F�Y߬��(f��@��x�bJ襜9�oT�\�Zw^��󧕔��::��Ǿ(������b�W����a�̀����Ġ��>Hj{�5+��RMTX�g���E� ����`OFK2�$�k 5��}���#��"HSL+�/D�{	s{N�9��eW?Աz}�D���d�8��r6�����X���	��fR��%�r�&l��C@q�%<��N�J����n�h���!�(���4���^�&�-���S|�v�E2:L�87��=01�wz2zDgj��D37WO~f٘��u���='�Q�@����Cb~�e��NjD��7���Pp�;L	��I¶�����b�]Дd��w��^p�����d�q�Ca�Ⱦ5��J�r)��iY<�-@���Z,`����<	�X�B��x������6���3�l��L�i�`e�E���=G���w@�䴓����n
�?5��j�V���QX���[`�huh	��@0��`�1��傭m��5G
cG�W�!]I�Ȁ�����Ї���4`��/���5����p��+���l*s�}�3��{��ջ]�Ta�?	�~�C��̖��Nf{���+Z��E�Rq�;S�wK���GwiK_��\�I<f*��딫/�끴a_/*�^�y��#�y����C���FP(���G,�.����Q��!s;$��z��<熆4'(��-N�3��(���b���fIC�gr��mu���ϻ�t�3S� ����>K��6jH|�&����́�����.�<'I]۵5��[kU�,n�'���#�ؘ� ^ڕ(��Ma0��?�;��������'l��=I���u��mTh��^:��\2y廿#���