XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{{��%��a ~��r.>�L�Sw]��N{��}�nŝ5�F�]��Ŗ�72Ξ$��6�=z�S���ޡ�&�nθ�H*�W�h�?��(�y��\Z%� �r���:��d$~�g�:��'�T4~<���I�_V�ʹ�f�<�qC��A�չ�1�V4�������7,_e��3&ŏ}v}ąI���G�y ���f��v�������J
��Z�*Q�����Of�e�QI�	^Kъ Z�s�b��<�I3��L�Qv�q#��B��X8��σ�����'f�`U�f�;��Pܦ�w�p��bX�,���$�U�K?u	�lb�{RD�+b$��!�)��
g�XĒ��r-!�3$j�gm&n],�_��a�&�N'�XJWxY�,�}e�v��t>�֮�Q����i�3�][k>raB�xO��Q���i�������G��K*���<����{�~���Oi��6i+�)cV���(Jv)����]T���D=� A�P!�ȱ^�@���>��NՔL>��'��L��) �yy��2Ĵ�Ma�����29��Z�G �` �u�2{��W�A5�@/�DÇFi����@\��kG�G�D8��v��jf��ĝP^^o������^�}('%˝T:^K���p�$�H�B ��'�.��r�Ae�f�(Z�2�@Vq��XY.`��:T��>+6Q���5���M2�9Ӷ���t`���� �Ŷk�!)d��d�_j�X������z�/�w��XlxVHYEB    78b6    1dc0Ãn�nv1�n}?[�ne�9X!�A�O��&FPD �����e�]� ����jC�T~�D�������T|���S�`U?HK�t�ݵJR8��@�Xq��o��@�j�&�)V%H�ٯD�ۄ/�O.�8y1�*�$�|%YD&��.P5JI�KKg���XZ)�;���^�V��p{$��B�*q;c>���\�j��@0�	p(����ې�?�(n=Ȗ
�V3ބ�xք�U��er�NX�l���wf�x����A`�G��T�� xe�T�J��'��f�}�~��쮦ٔH�����_Ad�"�������SV�]ᘀ���zeюS��I�},����b�qH��OU���W���;[�A/�E�C�M�<
�Ea�5ecT��ъ\e��6-6��K�E��MhTb�v��Z��ѹ�n�Jh�{�6:�4�"�q&�.�!�[���"i�"n��S����#ю��+Fk�^��Z������k�
O����L��ad!(��nL^��"m�f5	�ϝrJ^,�l������o�p����L�c}���䢅�m/����v��(j�e�,m�64������iMqo�~)r�f��9c�yP��i5�dX��/�Y����;�zڋE�;��v��$�0�/2S�E��v�Հ��o_+b�K:=�05��`qt���u�7�RP'��ۡ�B5{�Ż���>p��v%o!{��K'���	Pt$�n�o^�Ktrd"�k�:��7���cP��b�fc��<�&Q[,t(��J�u��9�o�`1�ԗ��G��ؼ���h������K[Ql_Z�������$�q�v��ʫ�=���E���������F�L����"fpK��uq�#�~�����M�I?%�7�����b�oIEl'}2(�k��=S���^�INm7��;%q~i��u\쿽�b����r�&L������I������w��������&�S�.�a��γ�j/�)��������4v�K©* 67��P��nA ��>L>rG�^��J����6���@+9YI���~髈5��B��u�s�5��H0����ݻ�,��2
\�_V,B}���e�~����h6}����>��*�5����޼�z�%����t�?�5q���n6��t���Dw���du~yZ���F��H�?ԗ�O	�\���OH3�`4=��� �u4oU
\����~"� �J�$��?��u:�ȑ,YQ_h�8X�]�+Az�U�l��A�)"��C����"�
{�wt��0ܙ��z��"Q;F�����-S�jI� p`����z݄&��Q�������
����|mR(*�:gW)��^�t��rY�<�tڑ�B[��z�Ѭ���N��JoP�2^F�f}0<�	�qN��G�=i���g��,H\�J�@v�u�5&�+��7uS� �%�nk�I�9J{���ŌPަ����2��t�ҍ�fP��e����Œ�q�[����dJ��ҧ�Ϙ?{�~srD�u�����i���^�gk51-���3�<bp�o0��]oV�;�PWo?��1Vl���/|t.Z��h�W�i�`�Q��}�e�`8��U��� ��l��0��ϟ;	}hN�3�M5e�|n�=�/Pp������Ͽ�7�����||��a�#�? ��3�	�q�%m��Ʌ� ����R�R�S��dر�q�!7G���t���Y¬VH���%h�G�Z��[R����iX��O�Y7b[�������*?府����N%YN�zk�*I�cP��(� u�o��
+S�\u:r��|�&�ـR/楍9���^�'Na�W����5�x�Cd/>�蘩��i��,��%�y�z���<��9���rӼ"�`���w:I���I�E��$��^�"e8�ܛ�j@�wl)MfI�|Mu�i&�.�LPK7d��&�)�)�[�� �����藢3�[�s�y�7V�up�O�_�`�% �|Ep�2 ��s������z��#��DE��&�B&�r�_��j%�g���!�{/8?���1�Suƻ�,+H��aIC~�q���
�����l9������f�0mA��b��V�wm��VlM��L ��4���v~�[�s}�<mZ��~�����MZ�"�R�s���� ��aL�ٶ�h��2�U =��Td��0Pj
���ruA)[��Ϊd۟��8).Meia��}$#ok�W��*�r�q��խŐn���5�6�"�`�v#�� F ���soj#w�� ����l��f�
]�lf��1���p`G\es)	�h����6t
�-2�|vf]_��APK�⇏
V��8��}QLN�G���"�������v[kE�n"�����X��O�²���5Isp�Ր
��]^�A�7��ۮ>)�r�$��f��չ4�Z�2�in]u��Q�tU�����dO�i���-�d�
��=�Rs5��">$��# |緐�,FB���v�i�1�}r$�X�k"�^�l�fL�h����'��׋NO:]�7���=�s+CV�䦫��#�¿��A��I��"ϋ��!��r��/�x?��3Yux���50b�����&XٵT{,(Q�ϕ��g�oj���9�J��G��k��iշ����l��	
nrӘ)N�6�޴y!�2��hG���ۅ� �|��0�4�YR��or�v�i��.�q��NSkG�&"���H�@������X�ܰ����)�n���)J*΋�5-1��>���7Y㕃�SUvLN��򪹒`�V�V����3�N߫hH�^�@&V��	��Z���������&��7LӉ��~"��`�ȯ\�����,�3K6gv���&��98N��ė�Lj��&WU�1!����i}�:�w[6�c^�2���{s~��rQ�V5;b���&��c},�5�4�F85
�ߙc���MbY&#͡ܜ�O)��ꖭ�,_7����@��Z�u�����#�dڅ��Y!��~����J�I���IF�mhc=��@��������Qp>#-'���S)��~����S)B�L�9�J�w[�Z��CR++�z����=�\y���l)��cA�a�����pwOe&�=��-a��8T�s'��:F�C��4�+�±I�Y���	�_�w^�]�=1�{��~f�f��sZ4%8�f���w����|Zˣ��zy�+E~�*V�-S���֨oFn[<g[���wΘ�Ɩ_f�4w����RB��R�VF�cs0âܔ�U�3��Lju���,�x(O%ܾR��o蜠NcJսơ.���d/��{����@��գ�\��JC��C�&3/�u����Z��Q0T���m�V4?����30���\2ـ��Tb��9#�g��T�����ҋrS3�"�ݕB��¡�a�aC�K���u�w�F��.)�=�G6�B�9�S���5]�[m��s�&̒Ȑ]��P��,h%��j�EgRp�q��&��З���n����4.�s0�7&���PKP�x�cўv�2,����86����l�\�Ip���[0�]��=�d�ױ�2QW���p2��s�V�(co�hx�ѿ��9-U�_{��7���c�"c�<�ak��=#k�u9r!B�ʓ~����'*/��jU^\x!�wc[��ڰ�}@5�!���!X��v��ZIO� �IYR�C=Q��u�&fVk�_��T��`n�p�"/��W��3<�ψJq~�+Z����Q�6�/Z����/�Rʓ�5�5�_\ "�`���'���w `<�Y���/�g�m�XbPL�����Z�s��_N�?)JR��{Xz2p� ��G����8�-{�l���3�5�������J?@;�]Cz�����L��c��@�u S(�x���ຩ7��d�G<`�z�q�����X�7��8�:S��r�3�x�d����:Ig:���a��� ݜ���{R�����;��H�(]��-#��MB(��6�f>��:Wx,��6����*� �n}�J,@Aj����g�]����I9!O�׫��DѢģ�[�?e�"�*KK��Scm��T�OGi\�Xhʁ0���l���Z?>n��EY/p�t ���<��߷�'9T����,S��⬨ܨ��8�r�-� �`N'Ű��䮊�;��W�Vf���^n�����ݥ����#��-�n�^�%�u8bo����67`�/�:�'	�S�y��I��-���.��If�
r��SDr^�>=W���8yF1H�vp��y���%�A=�є$el��=�M�]�ZG�y�H����Aѯ��>�r1\5��=�������I������F�řs���'z(�{�޲�H�yM��K��(d�Q�3pMφ:�
MX�\3�Wl"�7.Tjd^��w��!O�b�)�f-�F���%�k�	�r��3��)X�L~n���8��U8�@jIFSuq���5��@�u(#F���5��������d3�Lv�=���)H1� �Ɖ���	��B��9K�������[e�� ��(�Y���Z�_�Q	�a(1��>�'��"I�RL�-�4�dyg���7!������>�`���A+�&��8�g\�W���L���YvL��;��)1\� � ���N<���4�yV��U�Q��k�#�c�H�G��2�l�f&L�^�H��D��4�2�A1��f�kD��F����ab5[_���B�J���<��x���律��qM�p�.���)ߨ��7��
d��!`5i��zɿ�i��78q�<d��A��������_�u�֊Č�3��������n*&K��+_�%>�����-2��J��	�G�+ y������C*á~��rt\kc��&��	��SK��|m3�$/]q~���2x{{��h2=`H-��������H���d{��=��&-����Sp�(�>�JB�t;��%lb�F���s�.3+�8�0�W�z�N?��ID���	�+7ʠ/���C�C�˗�oeY�3���r�^�>�2k����TI�E��g��%�Q��!��Z�	���O�܋��F+�:ӆ*��&�`'�z�5=�k[�ky�H9�u�?�y�h�� Q;�^7H��G��[wE�D#�*����&O#.��qs��pT
-�"��@A?*�CS�Xm��&[d<?Skq��<�}.�P+S��0��q1�b(]aI2��	tE����i�2t�#?'���^�su��;ۛO1@i��Y,8F�KP])�bq�F��U{�o���)���Y�L���%^_�۽����x�	�v��.�6�~���y@������Ԏ�H��v*?��N�g�v`�(�Տ���3{o4�Q�:CK,/�lL�e񕇐���b{2= %�(�׹���9��i2��׾��5�h��L)����]IZ�rי?4�))�U�p�O'��$�ŪTc�V�?�KC��"��>}:�N�?��J�_�L�51���X����?H����MtW��A�/!ͳ;,,{y1��[��r|�^%�bK�m�C]�`^#��Jx����G�k���=u?�#�9��ȫ���Uw������%��y�m�:H�h^�ꌱ-�9o_H��mG$�`&��{��v��@@FR�Ut���Ш\���0?ن�R.H�:D�M�+��������wV9ݔѪZ5蔽�lj�@�Aۗh��%��ۿn� ��R��Q�0�	{g���rk��ikI"�δ��o�>��v+���D�%���,��;4��:2�k�GQG93��(��R��)�"C�b�p`�G*�4S5����e�}�k��y����$bO�.P��OR?,L!�IX���3js�#Q�}�Z+߀ť:��x=��J;X�Z;=���s�W���ԏ�NώG�Q_�ei����j	b̂ncc�f��g���α������E���(��4�\|3�{e\�����ǫʟ �!�zO�6�^ham;��"9���\�̵rg�vF`&����i��$�U 7F#��e��=~��ZƂ�D8#��aP�ֻ
�:k�"��^��"�~��c��ھt��.�։�m9��>��N��e!�4RlN�ض��H,8h����S�	�ܜ����?���7���C�(�|S?��Ḽ�͋*z>��j���N 4��������a�g�q�G��,��_��m�BR.Ss�}��B�n�vK��a0��}��4��I�aQe&���WAbm�����D��L_?)�i$'�7a���Z�{#
��;�o�r�:z��Wt��>͈Nˏε}��6�������3�G��c�Q}BΚ���� Z[���*;G뽝�IҲL�ď��1|ϼC$p�2X�7�tE.B�4�(�A`
��wͰ+��XC"�����e���A��L2L�7W^
b;��ww�-����hɉ�7*H�S�9I�?v��������~�FOڹ��@`ۼ��7�áT]Qn��Gk��Pi4`����T*K�)�WZ�\kY1"�XB}é#@�:��-��d�����yG�����8H��
}�h"9�p�c���Aw�Yl�������\/�QHW"Gdw��a>��&p����<Xi&b���3�{)g^�[�k�$R%�sm�k���2#�9��B��w��G�w�&��p�N��h�t�湫&���s���\�R,�7Z��� @����I�y���a��ssd�M���8�iK �X���~�{��,�^���H/����� 5\�}��4��P~	h3Տ���N�`�j$6�#���Čt�|������t���{zw�T)\�D��J�������M��g	����ݪx�L�z9w�޷5��{.&A|6j|qYF��#�O�Q�z�,.[�4+w��\�p���V��ʹ�yЅ�'�<�^_�r��G��ΥAϺp�4A
p���ZX{#���-�$���vF�be߄T����jG�R�Uϱ]J�r���^'I�����c�+������Ft�і���V���J�����O�L���{~�:��A�e�7���r��9:��l�U�f�zP�nv�D�$+Z䜸N:���%	��&0�XG/�zwW� ��ì{���sce?Q���;U럓 �Q �\8���@��e_��+	������J���5�U�x�Le?f�@�U�ͯ�FJ��A-�G?�!2�=`��^�K刿�T%����]'EEY�f �q<���RW��Ѓ���A a���.��� );�Q�`]�%�T���l��1۷X�����s[㻉���j���� ��e��3�}r�aN�y`�b��ẏB�GLU3y$Mncp)b���ʠ��?.� f����.�Wx�k�^�? ��?v�'.�����H$'�8=9��y�b�zl^|%��̳#�������f]Pε�����#+�,?�v��/���4��ʄqx�pK�oD�*��zS�W9�����Uj�Gv�!�	��K7d#;�����A�5�/�XyFt�0���ME� h��:����<D�����֧w�����.