XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+��&?8X�]���eBC�x�ٙ؉�����/#�~O*�P*�2���:d��pz���/Fq�i��)y�}oܧW�H60x���b�"	�5x�kR(��v�/q�NZ#�E4��e�3�U�.�	)7��r6�2�`��꼞�?Nu�WfX.G\4�V�x�2ې�f?#�XŞm>1zh���\,Z��5=��7�ڲ�K��"Ӭ�8O��K�y���t4="�e\�Rr6�ݐZ+�i]��i����I>Ac80�Ww�J�~�}�dF�4�*/!�l��b1=�8� �ӳ
�������r�\�_A������Ƚ�yW.h%�(�AV�nIP�g?�-��~�s�|{�y'�Ի^)���B�����a�d��;k#׋�s���-O�h\q2�@;0*�gM�¯?��#Ê��g�K�#D僭f=K�s�./�՝�I�'�ݟ�=�`]z�h\8et���HIa�%�p��3T��3Xzo����ɡ�i�hE��d1��ԥ�Їz��1��ש��xz�d�T��ۍ�uaPHi���f�����S��H8M�zzV,�6.��#]�)b��廿�U6�&��T���G�22&����w�~O7o��*o�֪�]{D��H��z�s&�Ui��54�T$��e,P���!���6��3�a�B�c����3]�}���`�K+���#��	;+�}R�`a����*`�n"�W�I��{
~O�H�m��}���d�����Ƌ]
�=�I�'��1��O�G�}��XlxVHYEB    8571    19206��t�IåF��P�F��d��j�:8�r����k��o<&'������d��l��i�x��>z�-m�p��Q��yU��[��<bSKzL��`���M�t�O2�[@B_��<N��lN	Rh��UI���3����Y�Vo�w׮ĕ�YW�e��9��e��~�8�ȇ&?"�/I�)ad��	x⧮A41�:ֵi�:>�7ZB��"���$�mw%�<!�W:p�vEvL��M8jh��t'�Fu�jes�ӓdm�H_�-�ز p��J�b�0a��u�'�iUtܒ:N�W)��8�7��3ƺB[�"�C+���׎<�A2�6�&����^߲4bo��_Z^/��P_����G�s�*�������p�i�4p�l�����������/?�<�F�Q7c���R�D���~�r��G�Gg$;�/���m�yP�eT�"6-{���X�"":l���ڤ�ۣ�+$ML�Tu���w}T����[�gs"<�!��'>��B_]�Xf��
�S#��M�Y'�<b��P_'*>b�S�ܽ����T�����R|�G�DW������Mő&���%Bv2d*�A�n}�4xn�Ȅ����y�E	A�5��բ�ym+���%n����In'?�&<����iO���9k����C����9��dt�d�[z=�NI2F���Q�8ja16�Ŵ�a4�����`	�����a�1�)�ƶ��. 0���U�a���ț��'�O�g.�!�t."(���˙t�<IU�%�P7{g�P��	���FС3���T�t�K��4����m"i�6�	a����?[dلw�x��h�`|_��j{@�tl�O�J�A��}��*A�0Nʭpbi�x��m�fW�1F{�����~fk�,��^�7��3f�֘p��#�&@ �(e���H�&rexͪ�ݥ-��:� �Zb�˔�զ!�^;nQ-`e����5�4�3)�id�$X�wZ}�&�3V-�\��Q�xh&:J��mx�1�>L}�TcH'q�s��%���H�x�?ir�!��~6���gΏ�W4��Tt���Ft�n*�\��veSߌ�uX �)�5�h���VY'8+6�?�@� �3�e;Wh%�p����D߮��q�p��ń������G�m�0�"Zj�N���kw�xʰ�ƞׅ #�PX�
IW˗_�hx��=��v�P�A����oF"�Y���Z���\���®Q5��y�3�K�N��tio�2� ���>$ڒ2G�3��Aɡ����dv��i5���h�Rϵ�p�绪� P�œ�N�꧐�[yZ�Ȃ�c��V�L���������g�亂�B0����s��'@'�Z��Z�N���V-Y­�YZ���<���J:��xa���S��&4�"���"�K	�|�q�:����F���/�Cx:���g�:�9_ׅ���D��C��ax�9k|��.�8���p׽�T�מ�J:�dAr�&y�g��f��c��sX�-9��Eҏ��l��LgIs����==�B�U�&����>E��ڎ�0m�M�(�r� {7s���[Rí\P��xV ���Wp��`�Z.{���:QQ`/�(�ܼ�:J�\��旾?��X��5����p��i�x�(m�(��/ڱV�vy���
_	�}�Rkd��"`�A��8��[�v��H��Z����΃3���@���q�n
��`H�n��{�Zkpܩ�Q�����y����e	n'�B�J��6:<��%�y۳��CB��u^�krj_S�2]��a"c4��N��@1����Ts������k�F�f�*�ҸWx�&�7՛�Q��l���*XL�ronm������n��)�(�[i�F���G�~��6��������^�%~Z�>S�'�t-0S4���r��*���/��*ڳ��`�Y��%z��m�FY���~���3G _��>��7ڀD�%��{��	����3��w'#GP��,���h�uGB�������=�QEj�d���׾���O��1�tbf�������t�,�+�79������!�e�BdC���S��{w��TA�D1j��:��h�\��\>(.Q�16gc�����m��>�����2�ŖK��>c���^�<���ɢ�s��h�Gf�{��
^��͆��F  d0&)�$�BPf��/����0���^�}"��HW@��>i
$��R����y��t��k�kn������^g�x���^���O$OZ����r��hk�O)�q*�r��Ƥ�߰�X��۾�Y�*ǹ[��)�.�=�?��O �-K���@�?�� V�M�d`V��o�!��9���ƭvv]I=��DA,���|��Jp�JM��X��
�������s�|��xC���>����|��<���B�i�S����gl��,VhăD�'�����eo���0EE��F����nzKu�?xl�\�F�����k� �O4K�٠���07�F����!�1c]<%my6G���1��u�܏l܈^��{t�ZxA͟�N��r�K�!��#���iy�|���臰���m�����^��"I��w�N��qc��L�C$��g�#2����t�@AaP%�fګ�f'~��B��R�L �"��8�N����ϧ\��Rݞ'�}�J��@��}��'���g><�~�����@�as�L?��--����A�,���)�"�`��J��P�~���kI+ �-4q�֠PA^��_�����@���z����٣�!g��[� ���_<E���O�ftok�2�7d�B/�d�"��蚩[o��B�s�a �#0B%�P��S�݌�6vV[�>��� I.V�fK��9n��� 8�uG+��Жq�:�bN��Rΐz��kDLNH���P��A�`A�8��O�'��.l�䩾� �zK"`R�=}�N�a���}K�������ƣ�� ����ߟ�vn|�\ #�n;��an�TT	�]��_Ʈl��`M�J���bIB/�I��l�h����}'OD�gƱ�>W���8�4�I�j�M�E����ř�C���`46N� G�ސ���i��yU��*���F���VP�Yof���Q���+���B;/D�ㆠkBlTh�ٱs�zĄg%o�m�T.�Np�*]���.�w�,ϧ��¦x!E�����t���z3D�'o��eb��e��g��KF?ˬ��$�^O� �'��P���*S!=[��|����Hn[rIj��eI~U��'{&}�E(q�I��8[ِ�t?�!,`X2[��(�zF��q�3��R��ty�<<q�fI;+�|�45���U2��#s���zC������l9Ӑw�3X$�I؄ HL�%R���O������	��f?*ʺz-�)KU}W!�����&W��'���ky���\��|U���&7��a��z�|CH��e��1([O������靌ڈ�J4C!.�	?�������q�6������%�1ӚA���3Ʀ��-3��؟�ϡI�?K�Ua�wK�.׉DTюe�Fa?�ݗ�T�}�rc�G�؍�Տ_b�~^^,W�o���l���� w,"�]�rk�t���_�<��N�i}]��6�k�ק��9f&Cw;�t�s�Z�+X^6̏;;$\�#ߛ(ݕҏw�)ٛ�1�uf�Rd��
ƂS�`�m�~��SPF������$a���6�	�F��E[�g*{�rB
���Ɏ^~kLR8H{�����Q�y��Y]F���_W�J���M��_:���8r�e�Oc��ue��#���87R��D��#"�Bک�{\r�����5>3��
+�����ȎF��L�\�Dv��Y緻��r��RE��P��r�9��H�]B@�BC�p�@`�qBO�A��8p���N���;~�'F���ڕk<��<��%mZS�����ؿ�\�Q��O���s˰�"m(ծ�P�l��ꂈUv����w<%��zB?ȱ��cK�U��E[_AUgϑ���׺۱;�mR��n?-�8���;�'�@"P9���	U�:�{�Aw�Ʊ���Ara)��=��Jb��~�^6	��2�]������Y��_Qn�o�
���}g�������iB�d����X���sڽ�I�5 ��O�7.j�!'���Y�?�'���6�a(�9����r_�M�d\�mp6������{7;)�q��E��w:*� �x��RS�����ԣ�B�c�e��sݿ�WN+$Vs�BvnQ��JM���I�?6������	d̝b�lx����%���(����qUŷ�k�/�wwj0��Q�V���ipX�t���,�����)�v?�O�pQw"�w�T�߅Y���t94F�P��Ii�P6EsO��h�(�����R�����0j�`"I���Y�5{h;����ԁ��~��u���e=�3�}��ڥpu�=[�W<>e)[���Vx�)O�ȸ�pl`v����kN��/@�\�A�"�z[E�����!o���,�����+u��� �#���%��
�2f�9���f����S��g;����L�P�ٗ*d�~.�aN�b��(V�#���nW�i�҇-������)49�L7K*OI�w�/ϫ��(2��Q��VZN�W�F�2�W��G'�=���P+���E��ܒ�\�dXm�ʔ����ߟ�N�!�v��'���J˥�Eh&Amp�sO#ct�^���Ӂk����3ic��Pռ�-ւ�Bwx@ʚ�w]��R�#��gҘ�{��>�r�|E}���<�,OAF��6y���Pt�UN@e�	���� ��]ㆎ��3{�S��(N×q}�8O��銢�3����T�&j�F�lK�5�$sv��@��CAo���p�_�h�N��7���Wv��g��4�AMh��	fz��\$*[��J�b/��D3 ��+�Ƃ 3x��Ƕf��K�V?url֭;��P&Adc�6�����O���1����:>`Q� �[߆h����@$V{�X(����D�pD������R[	��� e��Y���$)��\�>-��E��WIL�GO�>��r��|��cƥN��@é��$����Sy�t��e�R�Z���,G��B��Vٛ<WQ�5,g-�ޖF�g���9�.̊&�EZ ^�w��|���&=�ٱ��;}��A����������`�,�v��$;ԛ`�lq��uS�s|�@��}9x�,@�F=ra�[>ӥ _?�Ʋ�L�}�N^���<x:|?�_B9.��H�Ʀ��S�c��G/	ŜA�V���\ �\�'kw7F�p�qJ�S		H�a�^j �T��`i#�\'���[���e�/r���RLY����
[yF�;c��m\�Y[�wW�Q5�zs
N���=�!�a΋@A�yF��i]�t�܇4r���&�/s~��
s���$fCA��k�8N(�|o�����M�4�lb|M��5�W��(Z���١!���f��A�v�0`�d'���3Ȼ3�lm)5���0�F�B�͆�7��,�zɜf_� �Ϩa�Z9l&�6}E��SU*e�M/�<",�Jf���[��#iq+��M*	˺r��n�!V�[���Õ�%�h�&�
9�,�>�@S�s��b���A�I=)�8�%g��T���αax�S`���vݫ�>l+��0a�
�Z��}�d2Z���A=�{ i&��e_Vo(�|Ыø)�"Gg��)� V�$����XMCk��g��B^T��w&�����d5�Q�α��کbI�/|O�J1I0�Φ�w�l�8�� �������ґO�^�bi�.�_
��1~��0�!�˓~V�q�(쿳�W�_DB��6�d��Fs���v9;�¡8�Cp�g��ee�sܓv���C���[z
�1�=-��S��.fݍ�5c�d����J�ٳ��O�VI�)^��n�4�H�EI�$S��k�����[|��H�;���<n�?�_��c�F?t���\*�.B��(��]b���]:�q�c�Ìc8�j��C����q)2�`�~���j�j��xz߬��_6��8���.ȍS�-�t�A[���ĂG�nskv
y�"���z��z|�{	7\HcC���Y�掲�|�-��4�=�2�ٸ-�;����ӛlE/��6�,��U��4�4"���/�e��M�_�d+���z�b���p�P��ݗKp����	�A�a��;+~�P�����QՊ��xR�+V��C�3L�����IڍGFX��x^x�ݖ�ګwJ)�:9' X��K$�<7� SZx��$�
�P�LA(�Y�}���