XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;ii�Kl�WI�ю��3�ǆ�v�ms���s��C�B+>�.����Y
6ץޥ�Q��MQ�����XQ�F�S�:�	�x'?��p�� g���v�N�δ�ha�pj�Ь�$z`ceIv�M)�
t�Y!���T���R *�ʛ.�ǘi%੺IԀg8���k�/��(��%2>a���Ж�(�ѥN���|���k�4e��_�X��)�������v��GW�	� D�;���Ra%�ؐ�w�˔�S,������T�)���V@;�8R▐��	S8&��cJҞLV�8�'5���S���^���YY#6��e^z�gi���jj�I/���9�9̖ו�Z��������EJ��j��5�e{C�K"��|N�߃;(S��B�t��yH�̥L�-8�Po��hv��s ��	��`Q�J�@���ѷ�u-2���gh]��כp~�9ß�I+�&��\��F '��|��q��è�kٕ@���7aV���[BI��R�)xu6"|ȤF@y��?	�!,<�揎�~C�lQ�inn|��
� ���M>�]����N�'�����$|_E���r��<���ĪT`�3h�u�G�l%tD�3y��v�,�O�[]T+�ɤO%W��87��e^3ݾE�h��ٻzҡ�Ü>*���0Z-#ofڝ����Ӊ�߼�_�ڗ�}��N3i*~g�L��[��<x�m��_���W���g�/3Nnͧ
rm)�)�F�D]������Ar���,m.�zXlxVHYEB    1a04     940�O�0�廇���}��USӥ��:�+����`�Vtʙ�+�.[��o7�Ey:�A,���>%���| �=C]H�ŷ�Pf���	��A��;߈�`*��֫����2��T+�9q�����٬�.6�Z� ������J�"��H��/�6�K,Z��j�vԒXGk�B����W��3'��4�sc������m׼<�wW$�$8a��1����g�(�H�h���x�Y��E�����q�U%v�.�+X�	���F�Y�6���1�$�e�����cP��]V�<�7Q�U��՟e�O:�'�Jv|*x�@9���TU�D�A�i��i>s5Q�9���+]��"M�62��ͳϸ��{L�  �#mE�z荑s�m�}�bAec�7���0Kx^����A��g�kŻ%�@hٗ-�!�����K�6� QMp�a�+��gL��T�E|�t��X�/b��ǈ��3ɳ�m�B�^�jl.j��q��k��A��h� p��cn�1n�A=��k�h�����YE���*T{�$�8p +(k��yT4)�$n��3PV�5��.D/����K���V��{�.�uE�O�喛\8�͉�+��h#g�(36s�T/f�*�8��L��CQ)�������3�}S��q���<��ò�r�ꮱ@d���_��~Z�/�����̷7��T��j9(;09�_��)��d����=����N���bJ�̚��bɉmؼ�xY_���5��B�E������������&�?(�j)bk`�=��cI�C��G&�[�mV���aq��3����o���j�I�Nj�0���|�)(�]��c�ɪ�V!�}�F�J'_@i���a���a�4�����������Q���K�e�:�zƽ�o��lt8��h+ri(�s��f8��+�4j$�:[�p��3Xj�%;/`�Z��>&�]��h�
�|���q���l}�D,A
Eq:Q�]�rQ.���_s���AI�n����%T�����t��yC���N��Դ"���Fmo�K����5���3�k9��U��b-(�vѯ�@��
���w�7����><��c������[�A׆_�U6^�K���7R�yaD�C/K\�
��W�ʔ�YХ�:���<�8 x���ZR��񉆟K����]���c���u.�R:����i��W7^�/����s ꔗ-���nna胥X�F�����9&i��$�������`)n����Vv��h�|�0`��R����s���nj�'��㒌�7��zP]=����W�h˶b�Mg�o������Ki���0��.Y�M�0ݭ�韴��앫�Na?K��	%�wAu��(Ԝ�ؠ|h�>��c���^gX���s��l
��ıDHwg!�s����ώ�B`nU���<���V��{d���R��V�>�k֓��Qg��G`ʲR^H�T�PJ�ƾD��-�S�l��� 2�w幦v`��G���'��(Hl.3T��?��z�lQo��+�`�6i�4�lw,�f�;i|�X$�u��+�(x�3���dpkw�D�߻���B5Ex�������ނ]�ʟsPO�z��;d����-����h=y(��5���Js��h^�V�\�, �u9�5����<��)e�V�
��/:�����M0�weP�0���uWj�qVEWr7�럈7�%����aP*#Q�Mv�Pk��g��G}?mN�h��~�ZL����lX��-ߌGc���.Hs�:��W���v\�Bj�g͠.������5#iJ�x fi������%"�/��p�q0��Nұm��]�bJ�k�%��/�����5T�:�X�ҫ�F$���AҬ��S����D5��Tc �P٦�搷B�ݒg�d2F�A�%n��\�09̨�F1������ MHTt�����G����e���DZ�)�Ӌlv84��J���I��A�$|�2�w`m,���8���oh����hA���=��lląE��F�M���	�TN%JJ1;�膦*�D5`�o��$�.N 5�䞇��VΟ��Z@��©�+�h�f�`畑�X�F(o%�w�a��[5�sq�,&.�*�Ay�|��*cA;��P�t�4yI���r�*�N�<�3z'�xþC+b{���%���C���-J��=�pyGF=+�
_8]�C&f>A�4;3����}��RV#R���Z?f�I��	Z!�'2��į�9���G�B����B��'�ʱ��	9���uW%U膏���W�8]��%!NC��l�HM� 