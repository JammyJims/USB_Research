XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��a@�H4�u�\ouO��&�y.=�Sз���Mn���n�� �ڹ��{�i��O����^��n�ctݜ�h�M��5� ��\��`ڶ��E>x?�ԑ/Z�_����"�ijg��j�������?����4W�^�O/������Q��S� K�+�,���R���P�f0�q�I�|s|�Ţ�vN��:� ���X'����7~9Ƌ�yq%���1�՚�1=p���`	�IT%MBQy��M��*s-+Jt�J��:����T7�L���'�k˳�»c�'�KB�6�*z���ޱq'H�@��^j囒,�<;���L�)�+��'��O3��C�98�@eYS) 3��.4_��/{���s��YH:�����w'�:u�z������qu�|�߄T�f��d!����o~� H$ig�z@՜�^�W��ʥ����ϋ��)����Q�=��C1@���	.�v��7�'��tD�����I}����pۨ{�>��c
��a�Y���|�in�� ���jyk�y)��)Ԗ��FM���:�]5��"|.:����/�B4��<�{H�s5��ư��S��M�.���ɺ�)D���螺u�0©�`����䝘~i��8^�ѕ�5����Rt���)�E �������V���@���q�_�h:��|HTk"�\�O�~D���z�}J$�ޗ9�m�6��m��� 3/�mRX�"7�����c>ֆġΕ�"��-
��0�K�� ��)zCP;�XlxVHYEB    59ca    1640���
�H)����xi��Qt�W pm^�^h�̿Y�b��,��I�e&�&��S�o��E%W�pW���Y���eqqvZ̕�fa���xRL�^ǘ(��V�5���h��f-9���Dا�_a���q�P�Ξ�%zYd��}��K���SQ���1m%�'d�x�@����/�H[�q�f� ���{B��&7��NZ�"��P�cGS"𶜡�O!ˈ5F��L>�^��N�pe����u�/����b=,g�F]�_�n<�cX`�2�~�O.%���#6|��ѾXj���4�q��S�؅�e2N����VTB7�b��lQO�.�V�G1�4����c`U�3��<�q
��,���R|Rr���Zc B�2]g/T���N��T�T� �#�Z^Ῥ�^��=�#��8��h���c��<�����G�/�XӃG;�߉QW� ��E�Ɩ����[�__�)1/H�GO�*� G][��@���Eq����I�ǩ��E1�\�4�qls��U���*e1���K�/�R���P}јN'���_��f�Ks�v �V�M���]j�����i�/l��I9j.D�������CG�B�����?��?�,��<�Q��}��� n�|�1C��Ve�-d�d���m��X\4�;>��.�lbK�Ijb}�K$~9��~�je}�J-)f5gA�N�q1�f����g�ݵ��ը�b����Xt��S����;A�W�͞�)�E)�`"�u�AI����T��<G��!�Ep_��K��1�Lf���/�:(�����Tq�&�E��"��^�K��������5����s���Op�t֋���	:�WJ�e1��?�Y�ǜ�c��,��r�݄j*���[4g��x��i<��'���K[Z�F6�,ľp �	8ٴ�mR��`��$gK."�F:X�O����[����L�_5�t��|"�Y�l�s��+�T�@�П@ě���'�[Q<f��
!4��-�Ż,�H�Ě�%�)M�Wq̤Pf���5���Z�Bi�Q$��{�䜃4f�C�b�T=��S�im�7�L{��y4�[oϾ��62��|8a��Y�`��o�c�BVz�I�Ϟm7�KiR+��_�8�ՍY�A�cj1��4�h�@Q�p���A_u�r�حO`L/5�\�Cm'�� �=��6����2��p�|�vTz���ϝG
b�����i�nB�d��5�$�n���dhu� ��*�nB��z�ߏ�	 U��;g�j�Z�Ѧ�=7��*��>��d��Y�VzޅK�@�"R<�9Q-W���o��&���w�8*�[�z��oU�t�V��K�2L��M����+�np�� �8\d�U.�=~�:���r�Z]eP�n)�ǂ$ d�@�?=�<�����i��q����B�>�Ģ씔�(S��ܾ�$3,׋�I֚:R)�Fn3�ל_\_�8^-�؊C��b�@�h*�jٖ��?�V�;�3Ͼ�67=���Z��0�!�t�O2����L��T�D������_��6fBUB�l�Y(o,��R��ل�\� �jy��S.��p�?m�o^��k�9�4��}��y��a���Ͽ�p�
h �L�+�?�>xp�?��&)Xǿ�.b>�N#�?�P]����}��#H���ԅ&�l�d�O;�.}�G�i�"�3��O���#��^����u�N�Mڲw�d�{���_���غ��'�{dw��,�÷&`�+\Y:��Yc���6գ��$��I��Ȉ�B6�����u~��`��^j�z@c�1�C�Wx'hƤ���}p��.cd4��´6�˶���u�TZ?'I����j*���1�[����⣁e��70�U1k�����"46ͨ&[)?irM���CC�u�GE;�JP+cJ��y�4H����X ' �!�<��Vh|�>���r�%�-[�UT63�ȃ�.������KC`P'}��-G)�\]JI6tTn��텈��V�Hߏ�j�cV��>���o��袰;�!��$m'_�&9��$u���8/H���_F�L_�{�v�Px��w'E��� uyh�Y�J��g��+�h����H怫z�&'4[��������p��~�?�w*�� �ڞ�~���
�Tx�.����5��VE��@g�W�Ly)��uu��0�TKE��a?��x�{�Ȑ��ߐ���p���
0�l	�Vu~�q'�_w������m�C%�<���^?S1�L���ZG3�A��E0�Lz*��,0�x?���KTا��Ѥi�ۼ5��9����k�<�T%�@I��ς��@ �������5`H^FJSƭ��W���>�������}]`����&W����h7.����S�-s̙��
��z�Y�������>�9k����8À)�s[A@=�6A��V�,R�.�a�:���	����Ό[WǁwBj�ic�3�i����Jy�kyTY���Sy�ی`��(TV�	2��?!,e�)"�S��ڭD5��-����k���dƾ|�"�_N}R@�!�۳y94�B���vZ-���:�����$JR'�����\�=�8�Z�^�3�(�T�5bb$x��Z���p��V`���x�|K�a/�i�6w��65ɩ����@����Ú\�?Z�h����]��Z�>>�~��8�XX� �q}�(�Z�'Ž �=N�΄
^��J�ۑ큌ͯб�k�z"�rm����M�ȑH�Y�0:������zen����c�k�ĝ��a�@SO�H5�eCKG���3�3���I��A?1�ù�[�V�	�:���%W��&��s���`����!�e�Pz�Τ�� I�Cdn��o*tU�ًw���c~r*z[W�c��ϧkISu����-�0Qs�@���ܨ���}4#�o����]w%�#����P�S��Ԅ�=2�x}G\�aG�������V�բ"��聼���-"N�ҫ`�?� &S���T�Y�&xz�Yu&>������KS�l(���EԳ���R�ˀ��L"�BY�8Ё�#7}
q^���)"�wY����uE�9�m�H���9��w�|������TGA�0o9�P��m|��Ծ�^-$$�J�Ȏ���7��8f��E���_S��Ȍ�������o2u�Wap
-�A.��+�˖�b��e�
����k���X4��_q�y�"��~�S���f���ʇ/� � !�$C#�).���mT�x��F�x%'(���77�rw�DU��?)����^�8)��s�s�i�[�� 2wb�3�亥n[�"�Y2��[2�3��~˗'-���$����v3�K�O��aƨ&<aM�C*<�,e���4��KF�dE0����Ы�Io� ��3�_�=�%�qŔb�a�{6���^�e4BfW`'�G� h�/rx�F���k&�C�,u��4����\�x��������C-'W'���{m���@C�ޱ��WSa�.��;��n|�.X���~�ptg���A'������t�?�}C���ㄤ��5r���_Wvi'7�����X�J7�<$�'�QU�8�}/�j|n*��D�^���ˍ�D/��EIͳQ�jWj^!�B '��~�o���ka�
�*5<=�2"�������ͽmt"I懴�3O�p�T� ,�p
Q\�e�`â{8vm���j��C���r��ǫzݿ���v�Z@�O@B\�Q�B�U�|9���D"����~߳�f���Y«�QJ�홺����>�av�1��'��O옇[OW�W��^.�۽���0�S�`V%�8qoAX������p�}�V>��nqOvҒ>p�8��`d�ߘ�
���Ո��re�|���҉���i��!J SACM���%�?��/)O㌚%gH �,V/RG���I�v�?�w���1��_u���p�)�E^@Զ��:�|����q�_��+k^(����Uwr�YhSM��8V���Y�đh��&����#i�_l�Q��ψ����	E�g1�+��-���'N'�E�'�x�'WȓrW?�_RW�\�@ƽ72�����q�(zQ������B�_�\���%+��p��z�af�Gx� ,�]��ـR����d�/�ߋj��1��e��35A��c'�	\�����J�srz�k(Jh�z^�7v�S�A�'
�ؐ���k�I5���A߀�eP6!�n������G����]z.�QDV~�>L���퀁�l���r�(�~5k�0����L=�3�Su��@Z�y�!pӋI�
�n6�@,�(/�V��|K��: vQ�!4��Q�>�)/k$�C:x��^�M���I�B_�qY5�Iv�O��T�B?�ydk(Rq�Z(��n_ߜí\$������}�E]k��
3�LA��e�X��H�bń?�k����re��d5mf�'!�m���[��ᑱ���h�a��&xi���m��nJq��U-c?�� �!��W����#���w�p����I�	����s����̄�l����W��^y�(���̘�'Ui�f�$�p�T}FqP�N��3x�oCMW �쒹3i�7-C_ȋ�	�
���XQ����V�~l
!�����!#!�\:%f��Z�
�]v�Jt��$%��Ƿ�����3���<�4&�%��r�wW��t{�(��dz!���I����{��
Y�}7��Ɍ�8���t��V���ڛ�	d����Qw�X�Ț"��?:v�w7O7��[�5�4X��4�´nhV��?�?g5�6��JEoM�����kZ_W�Z8J��߷�C�T�jH�i?�Sg(�Ҭ����=�r�2�p������
��[�9.�?Ś��G`� ũ<�Q���6���I1Y��/��
��r��>��`��7�d(No�5�nbA��s5��벽^��9�P���c}̱���[BG�J�R)���eT�p��(#1'fq��)�k���ZΒHY<�cɆ
@�� �)l|'� �W�o����N�,�q%���q��P�_*���"��F�z�z�
���YD�q�K��#A����M�Ι�	2ĵ=�����me4�x*[�j �m�ㇻ�Kb��>����""��T��!>�a�Q�Z��F���Û7�7|��F"A��L�N<���|@ �VĖ@���5a��)����o�$'��X9���X<���C[Z"�ظ�U�������� �E�Ӑ�\��qj�N4|��X�,�qȰ�*EOt���t���嵦w��S5�������W���_�	�a^!Վ��X�܃�[G�P;�է ���?�ↁ{!�Ϙ�`�v-���߳�k/X-G�O68�(��#h���],��|�Ł�X����(y���mj�<s|f�SʾcDT@�w�}Uf�$ƳO0�?79sx,��V�.�^��4mK[Ϭ�Z:�?��."��dd�I_l���flg,��1)�u�X��?rdN�K=�<���P�:t�q7� W�"��t���i"0����/�$硣h[ۨ$���ӛ�2N{����M?�s�/��GJȕ��a��B�h��g~_*���a�D�F�X{z��-�v�O�h�b?�_&�����b^7U��0G
�