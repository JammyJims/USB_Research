XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^��d̺]uʘ۲��/[D5�|u�t�O�fI6��l�187�Zh�8�V�g�7�[�:%<�r��b"�� Q?���
��}!�Z��$���V� � -'ୖf*��Q�n=�-�NB�^�_���l���:�Y�J�˨ā��\9 �'�z��KjL�x!�޵R�No�����Y����.���Pf�'�����-��sԔ9����iĨ�2Z㇊R��\q���eq��x���D�Ҟ� *F�������O��(L��Cu=�A����
)� a&��zE��m��,�b�!�����h��xkjI ������,(Qv�ײ���L�UM$��w�~k�%Ճh�$0@7�J�.��L�|��n���x��U�Q-�Tl�.����DH��
Y�\�혦��AY���c?pU�D�N�M��<� q���-n ��9�'�.6�W�fT�����I�s��iA*�%&���xֺh��Q5�o%J���G���za�b-��W=%����h�qώ���Ѧ#19�#�NTvP���!��I��4��'��'�ua��5��c���CI����2���+y��Z�讶�[�%^�v	�4/,i���?R ��!�.6�l��׳�v�r�iC4.��.��d�wq��Q�����!������7�y�.>�3~��ާ9��7��N�xh�s�R�����_��ۼ�s��#Q��̝14����+���F�-����"+Ӈ�P���rey�k���/N�#�w�%���<XlxVHYEB    287c     d90>C{�p"q�K��<�lq
�L��N=4J�`G���Y:?���=��FD(9��꾎�y��Г�벝J��Ո�2������D��ש܃�3z�Mzp=}=2��������v���:�U~�Ԣ�����n�q�'YO�m�(#E�m(I$�e�˲� ��3�NA| J��eA���h��Z�E��{$��V�1%��1��������v^�?��Lvg���-n��� 3��j5�0j��̈}�J.�)l#v���o�e�g��+\����Z��۾�Q��</�mXt`��b�c�R
���v�����`Ƣ��טl�CP��������D���aR�rOߕ��^GG<X=���x*A���K�B��D�jr)M��۞y�q�q�=� ��~Cv�9��Bi�Pj ���s�G�
fݞ��|D�����%�OK���O�l8E�� ���փ��"bЎ���HF���(�Bo�� �cZ�Ti����rH�6|:� gH7,�s��szγs1Gٖ�D��eGy!�vc0�1�
<�q��\p��b�S�%��:y�G$��]9��'��*
�h�$���+��#��T��پ�&�N�[Cg�
�uڀV$�Or��:Z�Az�o����89C��)����TQ�pZ]x�������r��a�V0���ֻ���@���<�K6[�B?y�'/^��âw)ŏo�Q��%��U�DjRqq������= ��X��f"��m6���T*��7� ��UE�bo�+>�e� z}��dx�{&�U�D�	;rk+��:3��&	�6hy���?�|������ҫ�Ğ��k�5Wn�^D�e����6Js"�XW� �=�an�E��泠�H�g�}ٖ1�Z��~��`eIz�0�/���BO���:��wUoQ����|����R3�%�Ԧ�|�����8�B�2W�2���qPW�$�|y���Q�7��u��G8�g�Z��@�%!hO�/��5H�Dc��yB���Q��u��J:��d+��2xIđw�wR��%.|ɾ%¼��i�]����wd�v�/�W���\�k|U�5���r'W�*ʷ���~䬆ppI��8��܂GS�0���k�+g�Vq�pK��>���G�xx���,�QO͑YI��,UT$O�nn��W�'��Ϡ����	0�Ik?��zҠc�\T�W�>�I=\�`��>�e{ŸXNPLVE"�_)�J6�շ�|��T�pH�BM׋�|���"Z�X�6�4�[��	�lҽ�^� �b&�@����:����p�>�8�j�b���wM��8]�m�^��Ыt�B����LB:����]i��w�ncm �(��5��~�2n-�4}����b����Q!��EMI�HgA�/�	�K;�D�t�a��+�ԭ%fM�Y�@&me�5E����(Χ�E��W�W���]*�$+�BH���Qh���'ʱ�ֳ��UL���j�jJCUZu*_SR�d�����	�X'5��'Ej�Oy���&��XO���`�Rg|�ʘ��nDË���>~�D�f�������UB����6���4}�6��BU�EL�P@s����N���{)�*c6���/L��U
ؼ��<J�*#�Q��3�Ș��`�O�	v��"���%i2�]4.R���MZ�vkU��=��u>'j��B���"�|޳�t@ó]ji(|	\�D��:��s?=� M�f���4�e�9��jq��~��r�l�D�2�)�YYP�b��� ���Z�4TW�hͮ�o��Yߪ��nW�Gρ�gtc^��e���E,k.�U���J8���>�m�u���,UjR�|]��GFa�����+HO��b�Ô^	~U䁜a��M�ޣѻ)/��Z+�����EM&\M����4�[�'-)�r\����ԙl��N8�qX�zРJ���!Q�ˮm[��6��F�U��k���@�y-�i�j�t�CR�Ť�)�ҨI �}�Wu����7�A2.�b���We愠��=�0e���^hjB����w����1����=!�����!��V�I�OK��y���D�у��פ�`�d󇍶V$�"�Xx\D:Uz�p
�x���[��E���g���s�f%"���qTcP�o�3\�P�%_z1&�����
�82�wA[�<(��Ѫ��g�����SFՈ��?"�f�k�jǖ�]�����L!pG����wաQ���(��VeU�:=3���HV���p!̀
���PO���M��Z_Ȁ3�������G�4����}��[�4F���1�5�B"����4a>��a��ș�y�4��0���H�&�\�Nޙ��鯲Y��h074Cv\(�K��e,�BS�����W'b��#�M(�2S�N�k-��ɝ�DY4��kTi�ܿ울�0D���4K]ć��-�0���ҭ�Gh���	5u�p6'兣�~Ae�\��5$��u=���m[v8��!/����h�3�_$��-*�,�<IY"W뮄��G��JKW���@� ��W�����_٤827�
�� �	J�Y�мJ��r�Ѡ;���b��C[�\��x���)�v�Q���@[�#�K7���t%�kr��[8D��:������e��}s>���	 ���nNN���ŉ�[T�e�{~�E�o�i�p�D#�[rշ�J����ri��7F9#JhI$��e+��P���ŭ���N�ncdF���U�X]��O���)�qT�����i;�9�������[����ꭔ.���ǚ���:騷1�C���$��O����-��hU�B	�����t�A"�k��c}&P�4WZk����L/SR�/��ᐂ��Xo5ػk�ۼI2�VG�;<Tծ�)���l1O�Gj̙ �;c_7;z{Tg8
�Ό0���(�n���gjq4�� ��hW�0!vv�P<����e�:t5	Z��FWѨ#0�7��S��~�L��>\�N�$�P�d�n-)J�^��0�c[~��HTfR��},��;�#`��O�4�������zo�������(i�T���,�����j�T;e��ռMz��_J0ܝ�b�W����jr�=D>�4��	�\�H��� �mY�W�HɊ�����ƚW5�" �C����o�~m\0�D�q����%s�c�c߉����cuh(P�Ħ����nK=��Or��T������o5,/)H��S�0j\��mj<���b{���y���Ӽ��P'��C�Z��\��z���)��#��V$���GIR��E�i����"�����}/\��g��Mj�@IM���L	�Wk�`���-�O��ࠋ"<�u�Ρ=�@�����!��Q�0i0hԻ�S+9P�%�.�}Q�|���8w���-v���*ui�vm��.���e�b�蹺��0�A�E��í�э