XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������:���)���Hz�RK������]�}����ta�,)�$�+kx�Nj#�q�-
-�c�e���#���=��$�ơ�l&��<�w_�PweY�U�_���T~��Ϳ���W�E��T�	I���s:
�67�l})�5=�Px�/y�0�8�H0��p&4�h϶w1��4�JDqiV�>;�(~�xC�76M����e͒P�����v�M�,�X/��k|�H�Jk��� �Nl��*���'��ݽ�W>O�L;�B�5�Ϟ,�(p�ַYH0�B1*=����N�9N�d^wX��"{�����\�h�]�����J�;�l���vE|9��|�q��8#ű�
O���ρ�T���C�s��ـ\��"A�%�\�ȐV��� �ձ��)��-Aw�y<G��4ɼ��N�En]��Ʌ���X(�W�_G^ �M���w:�+s\��`�V�~�1�a�_G�S�z^�o|�1�%�Wlu�a��M�eu�4�����ׅ�7�@^�#Ԫ"�k��a��m-8S���>�[���K_D肗��m����q(����wa�}d�(�R�a�I�"U�����h7�С���<�{
ۓ�]�ltچH��>΅ˋ�d�#(�H:�A���C	���f
2K���Ǿ�-��)���Iɟ�'�8d�6"e�0����ڣ�݀����j�J3�x»��A�)S�#q���=��X��_�����v��(���LH6���Dv��lڐ�����XlxVHYEB    3525     b90m�$�{��h?Nuxn���;+�hg���4Mg��k��t<�q��
 un抜�:k~�X{�[�_�Z�6���#^��8��~�F�0�[jW�����ϗ�v�7�W��tO�V=\w#�^�F�� ���i;���49�
�Q�']���O��e (b�� X��p���-H&vo}2�H�3�_�CqB����'��}&'�ׅ�{.vQA��H+@��.�9�}@�l	~��O�9v�	 ���[-Ѥ`B���ζ�Wz���tL� 9����� ����	� �J����&K�S��e�Iu��Y�Ń3��A�^�Ð��D��^D�E�u�ݗf��~�Ro�k!�m���灷[����ú��z ���uCP/+�r#�
�\�6��C}i	QR���Ov���P^0Jߠm��U'}�pO�LjW0z�%9h�/�b���[��]�����z��q[ �6=[���t���q�hD�(�`P���9���M�P�Z������d��`��6T�$n��w*/Y� ��A�bi�L��� 6\��\�Q������b���F���k[^�ݾG���ϋ���	��W�fQL�T�h�
�� �����v��v�Q��b��r���ݫ^�?"7~���#GW�Q"�+6ө�$���KqS`	bM�C��<!5�C�pÄ���<��	���삢5�፾�^k5Ž|�ޡ]����Zj_�g$A��\���1�6����c�aW"��[n}<
�k�>n�l>�%��ҹؼ��>�9�_ڸS��D6R挏RGBY�ҟ�D�X�]���e�o��q��"��^+��͎�������J�?PH2B�%�$���X!T�(���g0��ڳH�,�w�h�SG?pX^��{���������,_����E��W�4SO>;Q�R���{�(�;kxlp�Þ�k�dIV�������b�csE��S�,tO�.٫�\ͮ0l�L5�T��,6\�ۗ�����l�J"f�L!�Bv�"�QSĊ��^�$Ȳ�EfôX�o��z̨-eް�m���Z'��tk,WGIo�(�K�����A�7y\K���b��I5T�@�D9��p���9)�=���!�#WT���R.�;VQ�u���y��{��.�?��*91{c�hǄ���\X+�qq��/��I~�*bNP�p�J^��mi���	��%���u�~>��[�Ż�OnD�g����>��؂���dTX ݲ��WlNgWP��N ��K��U��wu�l�S�>T�)#��tfAK5aw��SGlLrS�2��m����v7��#��D�֤Vw��L�Vm�� �����4�"�}3���û���UP�p���?Or�n��ʌ�i�A�U�R�|�{(��G�%sb|I�զ"��u@.jt�>������Z�"{t�y_����gP OF�w~1 #��Z?���G56�F�����o��ȴȟ��u)V��X
*�A�:e��Ez��
�'������&2A�� ��� ���I���^�����	PS/�0��q����tgM���B8F��H	/�;L->���	��p��ȥ(a�BR	�m��j�`�&v7���L�!$�O�Vl�O�ݓ�'B�Ԧ��x���?��+�D̕u��k�j�*������=�� IK���� tt�a��Č1l�I�n�i&�m �0�.�Y��g�����'��(����y�P�""�ҁ`�|�ՙ��pD,{l�7U���&�3�����jd��5&�9J`�D��E���%}>.ځX�T�U�¤
7�.a4������ə�c9I��B��V{���<I���6��}u��{��aR��W�po�̽|�k�,���#�N'��z�KɃ����yX65W�TZ�Ӿ�`rQ3i���Dl���T*��{qz`	���ֹm,6�<�&ߥ�Nf� KP+D�S�y�!L
�� ÑN�	�v�����I�n A1b}��G���AO>F���ZF��Ƹ�9q�ϫ���^�&>��|� :_�{��@��"���=� �O� 緜�����f��l\���3F��[�hj}^
��{� /f!��(�|O��g���M1�&��ޤ�B<�|��z��a���Af�Vh�8)ukŌ8�Y*�__u��� $TZ,���icj�ԱXZ�T^�"����L�(߈Wqo���ּ�вRp�ڣc�c>d�S�j8/�t�����߫5, !C]U�{���Z�׺]���bNk�����������ݢn1� �'�Y���V��R����tf_h�"'0�h|��?P���]Hxe�p�[�6.�F�xn�t��� �<P��D���k��م�����E��p��O�nxY����ȎQ�븪Ibi4|�#,<�s?��|�Ö�e]Z��Yr�8�d�v��h�FH���3����m.ıp,���7X�4���V�w`+᧰n�@#�LL�9���׍���@�%j���6��xIg�!��OӻѕV����":V��BC1��-��i�]���2S��-B�)�FB�VL��eZ$=Ѝ���	]N��S����@*©n��Kc�{��wÄT\�k�I1a3�����S�Q}�_�yS����)6�)�q�ԕ����d��$�X�w4����阙ff=�PZ���U�M����D�B&����Ԗ��tE�p�9��|���6ejhj׿�$���D�����B�/�^�4!�x���Ӵ�;�����r-��F��k���N-Lq��|��MDH���fS���6��Wlv�-"��t^���De�.��U��� ����Ž;'V)�o��J�ը���m������C�A���E��*��� �gE�+!�;J#���b�r���,H�\�=�&����P�uDt[h