XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C�RϚPn㕮�B���7�~��8��1 ���0�<��[�ב�ж�u�A�:���Y�
ǋC��r7�����_ê�����X�m�s�h19�#Y=�lo�>�S�Y��K��z
��CRH+�b�T��޾�P{�JڧdC���hrZ�A�%���x]���7��|}�Vc�L����^v��U(�CB���V�& ��u6[,�Ҵ7�r�Cř�\k�g҈x�YC�g3��� F�˜�V��ϒ�P��J{��{z��P�,�l�=N8f�����<��ey���#8X/0ߧ�*�^p�m�y���j���oz� ���;1�ѵ��`k�%ro^[vi��`��Rx�����*�d���|W��������i�S�%|��;�T����;52���I4w���W�r$+�$���͢�u
-Wc�wD󎖻�J;��8n���(�{��~��}ҿ#%t�<ѣ�8ػ8�k^TLr=M¡ךS��}��K��S���Ą�&i�������fXO�s50�P{�U�-u!�SwY��ϊ����z�G�߀��:�r���Dx��+PP
�}I�P��mxXN�/��͠���Rur�ڡ�6�.}�����7���s�D%�7�$���;{+P�YLo�����"�Ǵ�Ǣ�5�G�*�.�o�qڊ������
O4*)���
ŪB��'4z+B<���? /�ŷ����F�}���W��xp��ϙt�c[ڄ]�"�e��Y ��ѭ�2XlxVHYEB    23a8     8c0���)��F��7�0Cz�Ö6j�Ʃ�;�d�Ǻ��O�;[���!'�jaP�o(�R�T�s�S�������9Z������s����Jj��=�G���'��f��`���x�Z��p��M�S��A#�,T�m��W�乕�;f]u��S��#	��K,Y·��[��+�i���!(��`������w��B�������i��U�z�-c��[�����<^�@�e�)�~�����OP�c�^`ݦ��Rx(E/�����y���n��B�~ܘv�#��x�2��uX8�YJUA��~�|!%��{2����5���@"�<���ҏ�\�#�$cS:�5b�s��	VK�K�vSA#"� ZZ�3	;J�{���'�5O�x��dQuf�.�H�)⿤��#�R��E9�0�	@-�dS�{�λ�{l�|�w ��ų�:v@��Ls��	
AH�=��s�V7F Wɞ��vC��n�0g�1�#b�dН���עd9l���&<�ǰ�[N_4#��b���Lz��V����f-�����!L�R���^)_�6�!q�)�s����i��c,ŮA-�!Z����2��F�(�E�����jq�*u��Y��B:�W4���_�W����$�L�g���E��׭k�_�2%�����KYR� ����)�Y����K�"2�,����[�����L��F��ܾ�2�թt���9�ʓ�0�'��C��r��8�ox�<��:u���IJ��e��^z�Me-�:� t�U�����G~}�'_�ll+Y������" �U�P���G��))I�?)�j�D�Xa}�J�[���%밓4�
j���'�j���[/U�/����v���W��u�:܂�OL_Q��-����N_����5,�5�F� ��ه���&+��t���]�4g�_������+#�B�����AʂX����̅*��˭)o;F���E�ZW�B��Oyd^����f���ti�Z"�"UH"�������	eLL-&���U�o�&0�K�eq�6��}J�\*��έ5��9Qk0����}p@a�l�d�sS(��<��R�$5���G|����¬/��ox2�5f(�;��M�0b(�{UM������~YR$,��1�a?o�l��֟��γ��4�K�e�O�r>F1�I<�mTh�����BTwq�K���TT]̗LU�K+��L6�Gն�$�S�äm�����e��*]�ɡL�v��/P �4�k��t��������x?M�:f������*qx_}��dgs1����fm';9�To�	=4�X*�
0$>��� w��/ɞ�|4�Y�����<�����7w�5��a{V`��iu�FՌK�͒�ţQȊ��&6�
�z�I�+F��>E-�=�g��TK( +G��c �1�S�̀����"OkؼPQC��m���b��kgup�+mЧbCT���8����u&.���&�MϧBs"�P
J��o��{��c��z�z'=.��P�k6 �Cv	<?G3�3��𙮀L�_��u�L��Y~h��qrp�0�)�N�eJ�)6��X:%S�~L�B���雲�8v�#E����!�)ޒ��m)W��i*���������Y�*8e���YD�I�x��Ԓ{H(V4.)O�f�Ҟ��(p�*/t�� �}��-"r�������#FVC��������C���H����[O�H�$0���v	(O�y�M��c;e�
�?��v��e�\��E�,�|���A*׸0� �W��M�aVG��p�#)(�^t�'�K�z�*QV�jN���Ըh����]��dh�ϻ�{�L@w�3��V����u��O6]���]� .s�	�9jq�y1�%���\Q���5���΅٪5ԟ�d���cm�1�Kb�R�[��֖�ǚ6h��ũ)�Zg�R,�� q{��gD�"`��U��;�0��T�O����4��A�j\�{��F_�$`Կ?��N����f3����������gr�Y/��g���k��V�$��0���MC��6#
�2t�zP4���Ot`w��[�U֎���{x_B.q����+��`q<mA�e%���)���eG��z2��^���G��J�j��&���k	f!�����3��`�j�֞k-�q/����