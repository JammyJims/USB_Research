XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<3���nk���.�	=���&�&�gC�Y���ߡwd�7t?Tqd;aE�.�9��ڏ9t�W��P#�����i����恷�J]�ȠNu~��z��rq]�m���V��5j�6�S����y���]�܅��^��#��ˇ�!r�*+ �8k� �x=n�Æ=y}\?��5;a֩�d�����9�	9Dfˆ�[�EӾ˦z�vH���0�)�1��!H��E��Z~pq��W+e�������JsI0���~}�<:�x��G�x!����$Ty��,��p����ƥ��I���4��.P���.�{@~�i��kp[�5eːm�R3K;}Ԝ�:���n�Ā�)� �V~#�����Y<f$��WO���z�w�O�N��\��;LEe3"���d)�Ul�����	݁��?�Ͽ��%��y�g���CN�k�/^��LOч���S|�@o
S�>�|�����D,/������@����c��ȞT<�L-����C]�?qm�z��!�.s(��3C걙��e�ܞ���8~��+Q�z��<���ؘ�~�U��wk�wkՈ��vr�>B��I� ��toD"�T7?��>I�����s����@Ж��MO�^>}9�e��c%`/G�"���w�	
K��ZR]v?S�:�G������k����s���g�� +A�G�-�kD+4��F�h�T�e]5"�W�G�����%��Q�6:��������Kw�71K_W�a�XlxVHYEB    20b1     b10�@���"ձ�@������G
�X�\ٝ�;�J;~�I[�� �e�.FeR�㈑��V��7��l�O���~KS ��jۤ��`g���(�JR��g�&�Z�b�#�Y��MH�hZ���q0%N�ŀ��c�Āq�34�e�U�>e�>.X8f�z%���L4]�Nx�QU���25�Ȧ�~W��
Vdw��p{��M#�J%�cJa�jY�2�%H�$�NI� �`?�u�J8+hO珎Z�����84��1^9h��Qw(�L���P�A@��
j�X��W!!��G�=�������/�P%V�p- u^k�s���|��~��$=D�KT���z-��+�dY�����KQ�:^vR��>����!Jo���T*��0�S>�ѻZ^�
�ȝ���=\O�[ڙ�}��Z�<N6�-������� �+�./T=���n�1�E��:KH��x,�Zey�b�4S�`��wO+fo���]�'���¯}"Ҙ�'�x�|�_�����f��.�.co��]��=E�ͷ�����*!�o�ƴ�O_%��	3�6�3��|�64E3�o���2'�8��*�R����ts�v�����N�Zq�3^{�S1�ZF�+�-������'�E/VM�o��@O`�����!9��_�E� ������4j���YI<�f���H����F4C}��^P�$g�3p�8�
0��/(���O智E�83��ۅ�O���T�-4t(�����0��/E���u(�)C��i�m_�]��6yV�����̴Q(CcoI4��$s�FW*9�XĔmU���`ʑ�B��}�:`n2C3�}�|1k� ĩ��HC�u�
`��+�S9����Ȏ����ԠW%r4������G���6[zy��l������61I��B���ɇ=W����5�pҖwͮ�����AmS�y�ˇI�'����{���0�;��.鐧�@����`·�Q���3�8IM~t�irC ��nM^�(ӴS�7��8!�[nD�cp��YM��_Y�#�+��_��+~IK�<��C��w{��f���������R^+�h�C�]ފ�y+p�%u��&�\�Tޒ#*���n$w�3[�2���ω�GjiF�T�ԏ �w�K����@������Įz娸@K��(�'#%���6�M�@=9g�/����s����$muvw���.��0t��֮����7JE��?V�x���ɂsOj�b����������{T괼����>�A���;W(ba�~A&�_��6�݀%��ü����OP�}�� 2�@+ `�֜��uK*��f�g��S>Ec��ݸ���Sܫ>�u6��6����P$�I��nc#b@11�x�6�y�t��n
|��6�h��Y����2��� ��Kڠ<�'���P�RA���	��Y��6<	�E�چ��"��B;��[���#nཪ}`�Ҡ�q�?vV�����R�i+��Sy.��W#j�ܨ 8']{y߯ڛ��ۺ2�ֺ��+� ��-���d��ل��*X��v�DQ+Bw�	�][�(@k<�N'�u|G+$��P@��)3�����Y�zݴ��C/o7�.����a�Rd�1$�$�����yms�9o2�F̗���^��6�Ѯ,i��xtb͈�Ģ��jm�J��|�BW�:��<��Z�/��,��������l��`����9F�<i5ġ�q:�5ݬ^�6�`K��9��^����/3��S&bHE�it۫��oDθ����j2i��6n�R�G2�ܥ��_�7��+�Nk�F�h�jHlT��0����h����wt��_J�g���Z^;i�Kj-�b�f���F�%=YZ���Pq �6$]߹v}��N� �l�������;D0� k#������j��J]�L*�6�:w�XQFqJR	{((j[�P���Tޑ�e��c.8<M�JV�p	 � �^���y��C$���Ʀ���ͬ��x�-��u2r37<]�!��?*�ҩЁ����>�oY��P>"1
��� �؋vĖ��MIk}�T1D��v�Q�5E "���� G8��`��{T�7A�K�R�� �/wWmo*X��8�	�~��󨟆k���� ���􎞴�'h��JڥC���)�\�B����.�I�1�� �YεX����\[,ǀT����\r�a"��]�i�}� ��\;�#(�:�\�c�q?/\��5i�Vh���)��PEJ��s����rvM�%������m�r��M�|PԬ��V� s����ˑx�E�=�;2t��6Z��U������B^Cj�'9�/�ūHc�	�,c�Ʌ'�{�����W��t�@]�@АU�|I���l�2V���Wǘ������pb����k$��ִ��diCO��,j�eFᚶ����t���Rd�ϓe�`5���䒳軩�/�S�.�_4��!H����x�sY�á���*R.�kB��)
1;�k�˿��[��ڑ��g��!G��aB à���T��F�5]0�}lx�ȷ>�a{ާ
���(�
w����c_/���Z��h/?�cĵ��˗wm+�x�D?�ʵh\�D� ��{��7�\���w%�ah��B��4��-��ﻷ5��詻%Ԡ�Hz1r��� �Vi5�c4��L%r_`�!�����1U<^�F%f)���׷O�gc��Q!�����|*�Q��Y�(������� �
/���B,� ���/5��';��CS��F�WM����FBS�E)�� 뷲©[�w��q�h��
�����"�������HH��\͐�