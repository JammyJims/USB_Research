XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��XP#<�;Q�	�}��v�ѳ�Դl��m����];$��`�gm��bN�r�"6��+u�%E����`��#0\���+m�.���w��,A��3!��ѱ�|�����P���E.��n�#?E�%h��U��x
�n!�e�g2�.Z��{���o�]�l&i�ȝ>Ez���(�µƘ�s�|��u��'�%��xx���tPGD�D��e�	�m:�1!�^�œ�:�h0����Y^�rt��l�c�ۗ0
�,�xލ���"�`86�R��s�i���\�e�,>���T�b�8���ڽ#�O�˒�����>�Q^FM�Pj������t�j�{�'#��U|����GPO(RC�.خSK\�;���k�j0��
S���#��=h�T�׼������o)�)�|8�F�y��Gy%����@+���/�ƈ
)f�}���1 ��B�Ϭ|]��|"�|m+u�|n䁤�
K�O��h0)E��H� ��,�Ȳt˨�|�L7�y�C��Ù���P�=����1��	������/�GM�Zx�0k�7��f�w���;��+U}��<�����M����O&�2��Z)� �ʍZPI�������F�	��3�[P��UB�l���/�#�OLBr��f����؊�[���/._��z� ��#�zz�/�ؿ>�LЎ0' ���={���R��1~1@*�̊Ct��OI�b�O������`�,��p*j�Z��e��]��s��4uE��lĺXlxVHYEB    50b2    1560��>d�@���r�a��@���o�HK�.�h_�zNeg���)���q/���WJ ͖b��k�k��h����?��+����f�F����*0�#�Ԁ	������ڶL�xL�vU[�lZ�Y��Zh�J��#>�O�C�٦�p��z0@��ow�E����u�B@]�H�L�H\��-�VG���C���>�O�eW@��m��o�"�;Giբ0����
\��y�r=P���)g&wE;c��<]d�$=W_Μ���S3���
=#�G�1�Y�ӡ�$_�QDCl"b�S�l��֭�4�¦?R��$d�@,��%��4����t��^J��܄�,4�6��t�n��B���G}�_T>��h��닯6��T�a��2J�~1n�q)R��� #������"ܥX��3x�P��H,kRe:����t��.��m���ٻb ��m�'9i/�k�it0�����5�o�&rӇC��,����J��;��i"_$���Ջb�WU���@��^^2�MO�}�vm�Nx�����!#!�?M^���J�!�	mW�,�����lR��˅tF���2�D��19����x�k����#G~��A}��qΝ_6�u�y��/�B�(�&���4]�)!*�V+(3�`#)m�Bw�*�v�o�O/��I��Q�Y�y��qM�ڟz�L|�c���bN�v~7��'&��ةk�-0Qk
b�x��?��[�%ȯG��u��M]䮎��T��`x�Ve������L<d�]���ߩ�$�K��&���u�����M�������2�gK�gd�Z�˩ϝ�P,Z�9�����<Q=���V!Zu�{�g\Q*X�c��`'C7q�vu�VL�����M�dD�8+v�(�;	�h%
�XI�� �ӟz���2$mo�H�tn}S�;�#W��F6�����:��'e�����O��_[*�Oi�ۮ����2S!�v���I,:~~D#fV�N�������V�����r'E�f�>!m�W�k�B�T��G��}*P������6�F{5LJk�g@B=�k��$��7�����фߎ���J��@��2�l��/�Ga���YT�dn�Ͷ��%]��G�wTm�B��.���	-ʤ��T��&�z\����)Z���cr��cHw�q��Л��{k�@���	����a��O�e���֤����ZfѬwN!�`N~�Ǝ~%?�����9	(A�`�g򖗸?�{㕝Zm�V��'j#ʱa�}�Ll�d�"YAM����,\c�M�� w�V�#�|r���ȝ��6v��R}�)+ne�������h���f��ì\����F�w{�P��s�ඏ^�J�꡿յ�VM���,��������U�V:�ǃ�NC���{s�\B���;,��7�GH�t��cl~'�j(kv�d����v{e��UY�o:]�΁�&� e�Qmn�;�>A.���x���t�w�%$:������#�nVNvG�'�
�CB�Cr`z}�-+J�]��{VV�FK���lx)��fƇ:S-��"����נQTo!�a;V9#FP�l��"f��;
���;���.�
�rX����ҫ_'����~�h?����u���LMRrz	^�F1*�l���O�Lk\a��n���?@��J<�y����'����W��7	hw�V&<G;袹��Z0)��0��%�%��t�xq��E������N�v��a�XCy 碲_�a��Q�`� ��ٞR[�'�Le�'�|�(F���gA��� j�K��"��X�vJ��������w{N�Fo���uvP-j�f������B	7��ϡ���~���b�_7q�4Z{����u��-�I�ʤ�|���6���IQE�_W��G�>�FN}R��wc��D�	hC #re��Gdd
��#Z��[��K�-V�4���+Y���J�ʇ�+
A ��m�~_s�u�2u�g��E�&S��:�iG/
���@��߉�h�)o�\���Y�Y�_.0�5��'��_��,p�٧�+����}:R[Q5��`BƇ6�PS��%��O �9u۬']n*�5g�X+�����_֒0P7�p���r��@X)�����<�UG�o��R,wZ��]qD�6�&b)ǁֹ���ѷƩş�ͦ7���ǒ�r�r��N�a��j��xd���V-�(K̞�:ȴ�+�r�^���m��.|fK2�N#�T�j|qT-�]��Ǉ�����b�Hʹ�"��4�s�&�n���ӎ4v��>t��3��F��2�2���uᐷδ�H�Y�4[U���h���U�$�7����E��p@wn��ɀ��Q3iD,����0��'�Xp׼x����K�м��(��\W.��&3�15�޼�<CK�>���7n?��A?=�P�*R6\��r�#�q�9X��=�A��@�V3�C �!A$σ���:��<�j:
�a�1X*��e�J9�h&<��or��e��[�bag_����Y<ݱ7Ly�r�����S�w/����J�_,��u����:�X�#�ը4n�Z;��8�!s=����ƶ�E~�����F�>��6�g5���܂I	#�I2����l����\�.CU�	�F���]������6�M��$�'(�{I\�H�AX�CV�0ߓ�X�yU���㺹 ��U~�U�{]3
�k�7r�	�㭉���H�LQZR�ڴ��
z:�����hl.�Y!I��׊t0�/����گ�9���rL��ֆ��^�o.�U<��S��� "�D?EC1��2Ht$e����?d�A��4���;5�KpKz�$˟f��J�j��IJE�ו[{��t|]��=$�_�l�pH�C��k�%��Z�1��_�c
"��5e4;�~�8�����F�9�##��4m��fOG���xxn˪56�%���:�u�Vhls?0r�/D�p6Ȑ����a,��9q���oc�B)s^2ZY����bA:+"����M�|��D4�L�	�s�)��, ������6�;�/^A�#	�&!�O�Y!6�Иm��Ԋ�������VS*^��~��҉�o�l���7g�ʭ����Ci��S�j[�\;�Vo���}!�<4��vC��]�t�T�j	j����BrF��0aS�'��j�@'4oB�z��R�5��$�p���r�zyd
8Βa��
}G��kF)�W��\�;��J��U�6l�������x�3k��Z�
�xͲ;���	��yH\s/ؑ��7Qq�c�R=��tM�B��fs;�a61�Y���� {hQz�XS�ef��0g�sl�n,��o-flC[�^�n��k�^,}�:���vc�į��Jd���N�^/:���G�Vr	�O�sw��h=rr�ILPD;�ގ��: Yq��&:��V�C�/f� ��[qT��U�n�v��ehP�c;�y�B
	�o48BZ�����x�nlm�����D(�*�m��e�b�x��C<������1%�YL1���^���a���yhQ{Aʥ������\���ZʖP��R7�b`��2�����i�!i�ب�]t&3!���X���Ȅ��� c?�k����`���T` �4X����U���n�u�.^ℤ��u6���s��`(S�j�ݶ4�Yߛ̠�8W�M�ql���\a_����dW#{MgUE!͒��&+�������Mx���,X ��r��V*��S3L��TcVu3f� ӣO�>���:���V��8�X��Q4f�R�	�����|/����#U�g�V�+�fZFS��w;]�Q��n5�ϐnv�z��\�H�»�����z��x�;�Gyl����MEs�h��ƩZ�hn�,�r�Ă��5��`�V�p ��A=,�sC��'�*���
���`0�s�d�ٖ� �0"�� ,�"��{m�o��;f��,J�<j�/�sb�L@��lu�}�q����BʉEȗ�_����>N�{����5[�3q�����~uT.��d�3ό �;�')�:'�g�����#���Qt����1颐t���	������:��-�Rw>���W1�։�v�U�������QpQvX�5��9�-���fY�i`AE.��?�xOP��" �wiี����o?��P�����=�?r�ctn��̳J�ťs譇��πԧ���:�B�d�0�?k�z@���[Ţpx���dx�"��Z���O��J��T�]~/�Uj �W"'Q��)^-)�NR)��b�Dr�M��:V�9Q�����@�,��-o$���ל`�7;}z=ԯF�����D
(,��~<_�*v1�2��u�Ol��M�_���6����
	�hOw��a�و_�� �� �,"��I]�:��C�kYS�,�e\�.X�D�U�X(B���sF���ђ��8��>� gcDkM�>���!����F���
��٤	�M����
T����[���¶� nx���~�����v�M���{��z�/O�R>v�lzۊ�� ɨ]b������E�'d�9�9�83�y��x��l��Լ����*Wq̆N��KS19Q-���fOx�+g�/vQ)�����.��<�%���AteJ{����u�@˗��_<}%�;!�r�l��t�^��Ц0��f�����=���w���o���^�n�Eŕ�"ԀOm|u�@� ���;��m!�H^: �&�Lx&�y�!�l@��5�$lL��� ��~��)(e�ڧ��o�&x�56�m����jh�v9�T�!�Ӣ�V�k�g�G�Dyo�2�-#%�A|�|gȣ�;��`{�^#�JkF�\Ū��i�J�܆�����m�% ���i��6�e��j'���s2��Ry�c�$�q��8��ݚ���
�����#����+c�(Ǘ��]��"{�o9dJ�QzdO��r��E�c���rs�%+l��-�R3R���b��jY�o0(:�X��`ڻ��A��Sp�vʓt�e;Ge�W�˴ ��h�%�z���]U&���
~_�`}a��_��27����̯��w����P6����ats�x.\��ĳBiұ�w �3À>1�D��:S��\��{'�����{�N�&o?��k�m_J���x��#0��-nJ�9W<͘�A�n�V�3��=��n��&%M��l���X��ʒ:�*��:�_����,��֎ ��F&aCҏÿ&>T���8�R.�ß���6-�0�\����o�$o��Ĭ�<27a� =U�<��`��Q��"����^+I獂��V@F�q�<�,��!x[J��Qa\ې��NP���<~�$N�qD֔˅�$u5�7���QT��8�Q&oG��̫�u؃�+mhЖ�E�E�5�