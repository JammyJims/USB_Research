XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������'��)\���>�>tp��h��9�n�q/�� k���9b)]%�Y��=,f�~�Q/�c��~l!������#����0�ֈ&v�Br�J�����߹����18���i���A�� �j@v1fӫ@�H;V�&@wOc�D�=��X��<Ε��,r�Po�۞�&���?y�j
��	 p0����C0�� 0W�jm�vr�w��&u����%�8�u	UL�]k]��[曙�;�j�ɨ���	M����˵N�l�	k���s��%��cyv6@��fU�y����b�
��T\�/�.z��;6��>}�V..sF9a���]��X鱈�����jG�*�mBV�+!�/��5����x.
HGl!L� �2��#҄D�,�eF�V1�4<�H�L9��ǅor�yGڳe�3��-y�Ǘ�H&�6�.�E�G[�R�s8m�d�Q����G� j��U%�/��X;��1nK��-��u�"Z�a>%�$B/^�� LM7V#hfw��H����$�v�s�MRL��i�%��|1Y��=�"����G0��ޮ�*��.?�Fv��g�4����ҏ�k��.gM�y�p`t�8pw���-���VXr��Y�EP��bo�5Ϙ��\����%#��QH��v7Y_�`Y�D��Ğ l`�y���"FY�b��>��v�p�$�%�gt�]L��:?���1�X�#�� ���UN��$��%���%*�TN%Mf���_\�1��o��}c�uqj[�H�=��%qx��)7E�JXlxVHYEB    1dd7     a50H3���>�-i��͝�����^���ES�}g���1ϋ|�?<DH��A����U�@�ѳR/]VUE��8�#�e�3iUz�pyX��i�$<.�w�^>㏃O���#29eZ�pk�m�_]ֵ�o-��;��l�Vxtj�>h��ؼ���:�T��_CB��)�C�$�A/�[s�5PP�:|���$W�G!��<�l���M�,�%�A�F6�E��k^�;�[)_C�8��tz�,��Q�²Qq<�8�8{������l
�-�]#-Ŝ�i-Te��or!/ܑ�x��9P.�z3�ʵJȈ/���X鐦d�ĴK�!�k�����`�𐉸�t?/!��8X�q�0\������X�$�{���ht4�1����%,���D�}�ioQ!�4*�YP�A'��t�#5O�j�t�3ߜ��~��i�Z�|��K�GmՇj��r��'�F��ȭ 
J����$"J�[Ra:���;&��N�� o��V������~��L������ۚ��;7qZ,���N�ߑ�~����S/RmOH6<�[+Ћ=�h|���jG���+z��qJ��!
V��_��\���{Q���wu��Y��2��핓ؒ��3�+���#��y����L��J�\�[.HWm�V�E��Qk�����F��F2�u�Bʄ��<�.o`�dgg����6�e�.��u޽�i�,c�#4X�s�3-t��]G{/�gig���9�)˶�[T�e���zs� ����mH��ٵa� �ud�y,��Ľ�_3�<��j%@;���]"�*��(���D��
YǏQvv�G4=:��o�:X�&�zO3�,N��9=�ָi��R��8Ifoͽ�����$���y��+՟�T��8�A<գ��/$
]��W
H���?�?�u��9,�Xq0�˅�hэ�U�'��6�*Gu���	�е�e!�����A6m���`2��V]�
 ����cm�� qjqZ���H���vR�-�?y�� ���e�ba�0ˠ�܁pp>��v�!�{Ë��X��u��hi�TfRC�WR��y_��Q���P��
�QX��.g~��_(/�	H�b\���Q@�my䆖/Y��i܃�q7@�.�������S�#oĘ�����p[��X؈����p FV4�w��*᪫�{';v�N���l��k���KѶ"$oRs[5�Hl��Կ֌��\�A(njl.�����E;�Qؙ�aOl��dK��lE� e�O�g��h ���甖�CW�T!��2o�(�u>)��~X,\���-��a�4��	� h�z&��#��^�Mc��iA�4�HhleB̾�T���- ݮB��Gez��]��9I����n!D�><���NU.A�&��V��=(��N2�&2u�]��GL"�"���NN
iyQ�U���|�٬���h7`i\և��U-�1�&�^͌�Z=v��d���Cڛ
�ӣ�/�4a�g���:����Ԝ=���Dŀ���f~�64�SnO* �b�^��ɟ�.��z�׌�Uj-`�J�`iF뻠	D���b��h}h��E���F@G-N�N���\nNe%=��U�.*�ng_�]�3�}��j�C���L��qԓ!�H׼��A) �ɸK���G1l���oT��zP�/uO�씿<�0�1��'�K�=G��8�}f�.�>���{��b�W�_o��%�w28�W�'HD��U6�Y�%�X���|Vr� ��F%!mP����r-�r�L.�>��&ý�sg��8�Z����=V��!4�jA�IϦ����������O'��|��V�-�	-��]��gI����
����j@�_V��a�'} e{��4��`�B �:��qS��Q_���g	�Ԛ�v����Y�1G>���Y�=2��k��w3�ZJ.Y.���V�j��%��"`�z��-�8368��(���OÓ��l��j�N,�H�����[7ۣj�ɠ�~�}���#�$�Ɓ�g�|rͥp�VX!y��:h��u��^#�L�E4��*���+�I��I~<�;m��:����V�%��3f~R��%i���L�5�ɏ�2�F��e����v|t����^}Jת'0z(�t���	$��6A ��J}�R?��x���X���$�V3�3��cZN�&o����%��&V�1�;V('�8@�lnE��O���kOE-��X9&:��(�6�峔f����c���H���Q��B�?R��K� �K
��v���6�ur8�nS����ٴ�u}"�oͺk"�a��fu=l�k�\-4�5�>�Dl��!e1��=�}{����t�B:(���Dr����zcjq�D�s�ش�Ѭ�kf����1�@�r�(9���󡱧��YQ�x�]4�L/�Ld�2��
2����������Ƭ��x�QV���j����:]�� fub�EݬE�*������H#�Bč9���F�Y�Hbk�-�8��-��jH2�[�/\��Tɐ�%H�1��4&b�2�@���&���>j�:1����j�9�e�	�OVi5p�Q���h��nX�db*��n�����|��۫��lx�K
x����Xo}q4$�.��X