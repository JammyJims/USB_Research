XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�=?�)�ɘm��SZ���>p�d_���)� �J\�!f�?�n�U"M~���P&>�:���O΢�ʮ|���n�C�D� M��}��ˉ�O��卺��nN͓:��^e�V9dy�MqK��u\MB�	!$�2�Vȣ�%� D�Mz^Gl�\�R��ND����Шy!;�6ŭ�z6v�R�߂��ɕ�_G��Q�6�)��27�ʂT��,S��Ej���0-�b���X�}p���\�tcg%�e��^m���K��{��tKIS��$
O�_e>�}�߃79T%+>)e��U{(Ƌ����ߙT�)�?�G\�/�����Ы���)��?��l"b�`�Z8�ȑ�aD�ē-K.%�\�Mp���2��gJ0��r�{�"��/�!�� ='GH����pF�".�rr'���~{Е3c0����6�0(!�@Yp#'d�Y�3]��@&=Aq"$l<z?��O�f� 3ⱱk�@7��s-5GK�����HH�D��N$��'Tɟ�ք��lpH��5ߣ��;���X���Ef�l:Lu+���._���H�j,�鯚f��ˀnA�>�d:
)[���&\����9���*c5��KHn{��h2[�Ӌ���Χ�g��PQ:���@[����|�y5</[�-�A��UK�]���J]"7Qc?
 ��q����N#�Zr�M��$�^�6�Fס�R/����!�c�y{�Z�ֳ1��ŭ5�C���&����la�;�đBl���}���XlxVHYEB    4e6d    1710ޯ�\�ޯ3<�\+b��0,*�]d或Q<��Y��oBq����h��D=���x\X�}tj��]ut+�Q�J@:}D��c�0��·�XRA	F�	�+Y�ۢ_��j���l9�~#]�\�]�"��䮓;ʨ�%����牨Gq��x �QE��(Y(LHG]^�I� BJk)�6��ŀ��8��1�#����;��a��
�q8N����]H�g֞�6�	r��{�03y���}p�A�@	o�u�֏� g�0�]z�D]5<�?(�r*�)Ր����|�N/�������$T�JWM�qL���'� W�ԗO����h�������#�����������t%s7%w�EBC�%���}a~�r��/��8uD�@vm^����+?�ޗ4 ��G�F?9m�&.<��C���s� E����R�s|ubV�\����������Һ�R���@���;\б����槢�R�Hf�]y�-�`a�T�5���iI�7���>3]4Eu�Þ��m�����\�Ku�@�~u��!�����Ė�+��i��??tA�C���K�aFU|���n$BM�H8[T�,U��?��;;MB���pfՍƂ�������n�;|0��[�}c�8�� [���Q<S߾7��,�Q`p�3F��z q�wd}9i�g������<���!�)��GD����):�WF� S��R#�N.�TQLP;���l5N�,��@d߭A�@<1�<YYC�'GAo U���Rr�.#���M3l�G)8�D*I�wx�*� ��{��M���f
q�)�L�n~Ot��_��ۏ�N!��6���b~�� �Q^j�VvgJ�y���]��������Ї�O+��
����� ��2��(���Z��U]��{�H5e���59X}l��;7��l4��0��	���ޅ��4ր��0�$��h9i������T\�'Y�|�D3j�Xj����� ��F�{L�����?#@��׫P E��j�:��7���$��v(� C�I���-�.|�~=�c�ó�i��+�}�&m	�?���#��t�q�<�K�p��|E�drgM��K;�X���� ����~�ڛ�u�\B�2�������/�?pǻ'�y^�e�R_�G��I�XR�yn{�{��d�01z�}��{_���+2;c�k[���f���8�J�r���}Q��Ɩ㩐�|��esJ��Qu���N��!��]o��Ǯ�B�yʕ� �������*_aӀ���B�ןO���\|V��K�t�OUV�e�I��v�H�3ؓ3�yO�t�9��l����뱶>9iw0Z��L����\`C��!�Jz�X�j���w��;/u�C�%�(�r�=v���9=g�tf��+M�׸RUM�%�/qg�y��h,�@`@�B��s�I����_�N����C�xۊ����K�hA�����:Ԃ�T0�x;�K�,�}�}f2qJY !����{�N��!{���JF�DX_ί�����>1��b7�ߎ�}��&��VK��5�_>�.���]��Y|����KAyͮ�s[N�3�&RN��c/����.F�p�Jt9�S�Pa���$Q��βR���J|��9�N�-&��Q0c�a�f��e%�e( M���ʴܚevb-�����T=�����	X΁��C�^�|q�4s��gR�����r@���"6K/	��۠�ц6�1�S6t����Y�-�8����Ԑ(�_V�6�7*��Z�F�[F��
�?��VOg�Ԏ�5�G���&�e12LB&���+=L��EW�&�B�-D|ѵ�(�����}����}�-��P�z��`�l�eKGj�È�XIW����},�x���Y����iڰ4J�}H2z����Yo>��¯� W7&i��}k����wRw�����P�^̭	��9���(�:��?�O܈x��+����l}�B�RJ�
�C�.���g��W�I�}f�����ѧė����6hM'̳�[��)��Tɣ�f���g^3�%N=S���{���I��ԉ׉��ڽ���eC؍'�@D�H�����0����X�: 4Y��n�ⷘ�A\щCI�/��}97"�u�f;���6��Y���&.9�d�R��l���I�l۪� �[��(��(�[�g��O��ҫ�߶}]EFmɠ��K6o�SuƥG�,�����a|��)�K ��Ҍ�)��G�z��Z�s��E��h6B��8������W۽U�6W�"}b�'J���y�#�x�W��:���}n�_�0S��d���`��GqE<?2����b���7�A�䈸��A��������C�9W����J?���h�H#�����P���V�(t|�׺�"�K�6C AY�G!h2�wgx�9n��*��������������[�x[ve�d'g�;^�^x��cץ����ėq�]���Ű\��ϵ~Q�_�1)�����M9�K�ѧr�oT�{� �/��q��)�""�d>eݥ��܀��|�c��\�_���s	�	�E����A}��{�x�\���C�.\�k�B��J��_Y.����S�SK!���C�d ~�%4ܲŲk�ܧ�a���?P�(N%�:DA�����]��wʭGVX�z.p�(e}���fO6�d���+��+�x��_��t���A�&�4�C
��e9��-������Ǐ��q��Xj�4����fh�+# �ݜ�Mg.�$n�8����¹V��U(7��=��.��s�+����e0���y�A�E�*ujG�ԫ�m�݇�R��,߄N�g%35USV�i�7uF�8@�Z_�dw��2���IZj�G>a��C��"%LV~:%�r� �&:��7�hh3 a�r�c��PD���#�dy���N�k^+��u�|��w�ہ��f,*Sk�<�7��-��g;[���EN�eD����n�v�1�L�/x&X!�3\�S��_��ge���Ю�0�H����6���a��c��>���jRҁ@��.�&PR���QY~Ok}ͦ���S����C( j��W��2�Il ��R��B3�Ow�x���"(����Z�h|���~PzF�'#z#� ���*w�!�j�,��ᬕ�ϯ�H���c����f$��G����ͮ��R����.����^Û���_�P��j�!״�ZQcXK�/땍j=`�4����Ua �!rV���dw���y�̚O�t�������X��dL�(.�D�W��0�#�>A�<�8�>ٵ8/cu��LC�>O�v�Q\G�[I�$�4dm\-�w����q��|[�vN=1鞇���E�z��W�:\sNL�NY0iop
���z�	=0dIM�	��I����c�o�Kӑ1��ű(z=v%��oZQ[�^�ۚ�Nx��9>w�m��J����e#ȤH��Ш�6"ػ�q�PT�e���v#��G��A@[�<��]�]3�i�1;�;36	�\^��ρ��ɑ���V�X����^9ͦ��)��[5B&�Y�0�M;鬱����i $<2�ix>�Е�n�DJ�X�� �~t�g��O�K�P꜔Ҟ�n�	�uc�!툚�	S58;'���o���bl����bag��0@�x �J�{�I L{�{�-�M�ӫ*B;Q�9؀���̷�T�2G� �:v5�-|:�&p5� \,l�^g�?�B�e����W�0����i��Wf��xe���:8Q�R�72�ۃ�*��S�V�dE[Oŋ.��>I�aǝ�J]�-s��"�ټ}�fCq.����x?�����q�4��Xue�y���3�	r��0X�W�:6�;!�]�g�:�|��푬�㐌���9c�k���M���0�=�lLc/8�$���Ep*��C�N$NV��]#>�������>�W�>5��d�`g��1X{����U�B�pr߃�E�u��"��4���yh؟�nٛҺ�ڡ��H	�<'�A�xn��J�e��3-����.���'㜌�Jُ����+�d0\̰*����<!A晓-�F��8��i�I�;�M�iS
��Z!I@�v�3[�l,g�]��X��>����5��/K��Rr�.ׂ���dr�$�◅^��j��$�D����}��d���zC�)u�Q�iǪs��`�Z�a����̿QI"���^����?����M��65V�>�WfZ�jp�ݳBS|ZV�ut���R5��BB�]iz7��K�JTb�:�LE���?���^�'4l�~ ��ȝ�ZQ������Z�[��;t��8��;>���2�D�|��qښA�8��D����=2p��؁�{g
�!��&<�YQ,�ƥqO�x��ׯ�x�����J�O�)��[Һ�`�ь�oԽ�t�vMF�=����@���ջ�dv%e
��˟��C��}Y%\�K�A�|VM�h[O�do�K��/� �dMb�N}����R�I��r��ħ+���.k��lq��~=o�����P��|�F���zy?�S�޼�N���j�� .�圽��Ag��]j4�X�Ԥe���7�]]*��,���9�F��G�w5Y��bYv�ޠ��5^*�u������I�mdz���WF]~�r�0�~p<ץ����w�����\`�PT_��ʴ���_�f�p�Y��	��gc�h�zOz�FzZZܧ�~>�{���R��_>N��j�~����m,���6o�|����cRƅ�o��d�Kv���ca��Ә�_�b)�:�+��T�m՛\c�������A�8���*����D,<+�kC���<kSꐓ���o
�@qځ��Xg��R��I�1'�B���"������O�/D&�����pH�+�(�]]r��j+���A@4��9�vd{DV���̨A���Z��5�Ѻ�Q)դi��J �!r�󈢵XG3�ᯅ�w�9����`�x��V�/�ʿ!1M��S"*�\ԝ�>�nR"Z	4� 2&����>m'��ڕ�� x�,�l3O�Ck3�����SP�pҚ�Y��AB��eB��h���8У�Kԯm�ȇp���0�mi@!/�Q�^i�9�m��������H��шQ���\q�,q�V[뀦!m߂Rk�NX�2\D/Җ
�ha�X�|��VBUx{�s'��U�k.��@N���Id/:��fb�
����n�n$zё	�!+���f�AkV4�o7���?f���s��;p>�<a��?ƻ�a00��Gɩ8;�,��s��6__��m��7�s���"3��I�պx�b����z�q���Z�T̍d�{��~T9�Ei���!��4oّ��ۯU�S2�k��������N\=��4�ׅZ^��#s�( ����G�`"4/��_r�b/{���NB�L�d=J7��ek��3y��A�Gy�6�۳����ͅ�k��e�Q�m��Y���|��u��u6�j���8��%eTuK6���_R�|���'�� t��{�,�ި{W�Qgf��8�X�Kq�[�<����F&��r���}��ʊcq�R���#9Q�y�.}_+�������.���5VpK!��L��g¨���'�e��kf��:���52�k
ΐW��/�E�6��&}-�P�B����A�`�=�4���L�"���a�;|V����ȸM=���V���Կ0�����0Zљ�Q8���{�X"PpY��:��p������ҏ�8����m����y}��r�5�9Cň�~9ͽo���3�