XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ��Y�d��oRȔj�*s���6�L�d��.�;?��V������H��������P�g�&�)Rg��(^�	���sk:r�U�v8���=�gB�=Y�zJ\��6�5����4��h��*�d)�~�M}2j@�%G=uj�j���l�����I3h�=��3��D�R���pK�J-7���uQ:����f@fȌ�����/z谹љ�X��̄��E��ӹBt6LX��C���Q-TxbtӇ�>&_��-{�c�`y��Ҭ.B8��i��M��g�4�*Z�W��/�>���m�m�En}���x��t"����M��\!}B�uF���,`&<��ä�B�,"�u+Ώ�<)ˆ��Z�-���>�IA�y�T��0Onњ��z�G4�Z$f��Y�onC��]p`ߊffN�؇e��~�G�g~A4b'K� 9g?k�9�ޏC����c�oR�_L�yІ��U�u.,OX]A�l��뭡��q����6��1���9��L�Ob>�k>!��y����g�MØ,\��8Ξ�\���[͋��&K���˓�j���F1�y�t�qn���q���n��&���Y�X�����6=���W"~��y�@Y�q�kU���g�|Iͼy�爓�o.u���~��ݦR' ���ۛg��62� B*U�����7��!N��
ө�>�s>,2:A�r��9�y�"��A
[���τ�o�]�OWk�ʳ�%<���.�9@!j �Y��ma�:���XlxVHYEB    3052     b80YёkjRr;l�ѨkWr�ϥ��im���o���9�F�R�WUטI-h��Z�g�=��Μo��������|&7sų��A{��N�i~Co+���Nr)o�|��Hn���+��ٓ�a��	Y��)&ިw��:=�Ʃf��KQU�gj�<ܩ?6��.�Oe�Ŝ(o�	�A��Uo�2~�ו����:Iq�ZbqZߢ�8!r�y���$�k�������7,��T4U3ֿ��wBE�����9��ga���7�v���{�ƻ-�6t/7{�8�7�q!^�d�.��!�y�eog�ƕ�~���uʱ�O|���z�ۭJ�Z�N?��H�݆�y/�2j���ã��i4��p�P�bǌ��.�ؘ;�`��ƞ"^>��*����<�ݴ��a�4HK1E��|��nP�v�����G�q�@!%�Ҧ���L �ђ�|�J\�4����jVmP��0�B�A1`Q5klX��:�Jf�:�ym��}޽Ej�{G�(1+��2�E������� 3��Q�6�����kJh<�jT�6�epd�PJ�ń+�A}�@g*t ���o��u]�����ܧ�EK	��m��'z�n�9�����?���21,16�]n?�uc�A��].���V�U�'J���K;�S���-�gG�k��[�_Bk�q�lOa��Z�L��p�[��U�.T)y������R��ٱ��vJc��B?��E�χ�6�E�w�S����>�y.������B�V\���hӿ=��l�܋#ǡ����),ub��������ڕ�EL��N�@p�y(�	c��Ұl���O�z3���Ĕ�wřVѓ�T�>U��y&�﨏<��c��?B���Qќٲ�<=�2�ǌxݴz�H84�ZL6�Hr���r�6Ϸ�\�fP�����@��iJ���H�m�}�)�:�X��)�S��Ir����is���V�4~=?��C� 5KDXf�˫�Y��5BNEit�vF����t'ΑV~Cf�e������ݜ���TbNv�fe�m���^�>�Q%E¶`+t�|��9�Ǫ�rp��QA�r����6���ͅS�"�3��/��Bzҳ��u���6��[sv@��m]�#ؗ�w��CF4�����������7�@�F�t�V��DG2@�QU��>���wږ�+'&��'�Ȭ�q�eyz��ɱ
Z8�]���Y.�ՙ*g�+ p�yI	���' ~�w��������+GJ��yq��)O+1�2���ZSl��ףg����Z�S/�a��E�6!��?���


�R�ŒC+�\���'�jzu@�S��f_m��t�k#����m��˚H%ݙ9�<�$��Eߟ=����ˈ���;ݦ�`D����7���(G:;Vui��r"��`@��ֆ!��4}�:��͝���hF�ᣡ�! ��O�'>�D��t~WY�������U�N0��5�ZM����>,N�{t��O�7�����m���x�8OSg����oa��X���U����<���: 7\)s9QMA(�n�����'����~�X��!,�x#�F͘������9�n,��џ?^�:��]�8���/Q;~�y>�P�6�J�;��A��w6����/b�>���E�j�Iq@~�<_]v���VK0{�@[���)s,ZV�-qr�`d0{�|#��V�Ш�fɛn��8T�͜O���ܘn%7�*��L���0�����t���hI��3Z/���L�Q��4ib���vD����h�h���9Lw�N��cy�<�]S1v�+~
���H=wŸ����/�5�*���F;�����A�ϊ�u�x� �A��u�ݤ������?����v*��Q�i�^� �\�AEh���*
a~++:&cn�#���6�C<�!���S��A?	I�>�>��
�&�7/�:���	Mf�|G���9q�C���E��ݡK�� �Ք�{NQ��lb`���8���0�Z�>�'BO��)����ߺ����>q7�7t�kk�
Z^���sD\\�<P���fD�v�YMW��;Z�x�Gu��71v�(��lEp����T�$�H�d���h4�4��5�T8�/"9��L�֡#]�����P��"��i��#^��0��[��B ϖl	��z�X�]�)�	��s�C��๹I͙/��p-�id8ʴ ����������Ogw��ݦ��ʖ��,	K��ݡB���K���j˶ڣ ۹D%%޹�j��=��4���{m�U��6���+ p�R�e�����m�:s�LS���;?�s�r�1Y�����sT�V��Ii`��o�nGδ����c��+����b���S��S{5e�^߲C�y�}�{�7�ߩ4�pYl(��5*��B�7w����T!Ru��|��S�K�|<��=��^�!���#k���Q	�m�Y�x�a殠4Ť�dI�<J`ҥ�4�G�e�L��D����~G3�űsώ�{6�hdD��H��!{�M2��ﲮ��N��#��ws�p���- r�0k�;���Ѩج�����|���%۰0�cs󚐚����1��َt2��M�u��(,<����\����-]����(�8�f�D]�ͤi��Ǘa��`��������{�\��#M��a6&������*k鑸1��:�����:�(ҋ0/�1��v��Ү�l�t�6��5Dvt������K�\��{FW��
L���Jl@B�N�/^~���Ì�:�&I��J��@�n����6��<=�ԏ}E&��b����e;m|�sY�k~vĢ���0�v�~8-0'��q�n��Q��\��Q=��TC1��b[B�({:) S�����l|5�r�;�D=؛\��J��MJa��Z̤������w����i!.I�^�