XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����e>��s�G;�lʜq�G�*��=�֪���?Tr���<YMD��g���@��=j<X�_��{�ҁ@��
[(���Dy(�d Sh��`6Y�b�f5�I��h�+��ָ���Ճ]�բ�S_�T��a� MB,$͘iI�Ȱr��i�P��H��8��Α���۷��{Ldc��D�9! �@��-�?��f7>�'I,��]�Ye}$�&}�䚲KW��YB������YZ&&�]`"�`n�?��#n���^Le���._�wt���%N/�Y���⧛��P�L������Sx�#�e��ʻ������h�pq���j85"�����y`oP}�)�>�<�xr�պr��1��u����'f�n�;vq>*:F��s_�cp���;RCB��aቹ�A����ц�G[�p��7�\�X�3;ū%��e��������3l��Q�|2�N�~K]D�l�����Op�����{
���a}*��+��b�3�o���uj?��
�S�i��$ ���L���J1 ��N�zZ&:(Y��Ѹ|��=&�}�.E�۟/�:F��$�)��K��]!���£q	�m���Z�y��!&��Z|15Xߥt�=�'��8֔��hg�����]����|M[t�!\�}=��z��6�.�V�JI����]ţg��t���dF����
Ut����E�,��E����6�;s��kz�d�	�S�4����㌭�XlxVHYEB    28be     9f0D����sۚ����hz��:*�s��3���c�.d�Ҳ;p��A��gU�hG�K0?<+�Z�AM1ӻÔ��j���6Y�O1���BD����<�i6�>�x�%q
�4�B�L�QJ"FN�7�m9��`�2��o�d6��u<~���W>����`9B�ʒd�%w!�$Vا~���|���!}劐`~ׅr �o���C��,|3j=-��=�~���Z�pϠB:�,�*_2�6�0JZ�YP1$H�3ya�b�f��Ì�/�����tr�#�v48m��,Y�r��5a��p_��[��2�y���D�%Zͦc�g�!�҄��)���ޣ�I�/��� �z]9@y?���ڠ�����Um��I+vV	9�#� �rޣ2!�U��2]������١���	=�����8Jn`c�dÈ�!���\R4`�p̣� ��!lH d����}�w�x}t��ި^
�~K 0d(яX!�z�����g���KF�y�y�Q�(G�eВ��¶俼�����87Y2��8=f	�H%��Ղ$Ot(�HD����_��Ur�g�U�L��J���-�0��~�!��[�����-M�$B,��E�)�ѭ}�q�v�����(�l`�T��7�-��p�4�$�H:�b���q���;P�s��_�1����8W1��-�O=�>�0�CR�AF��H����}�����t�HH��j�F}px��Y�,O4��R�).%x։ò�D`�=����~ޞ��Q��LYޯ��<)=�OvY����t�~4���.Ht�)�p�U�*�?�rw�y���aװR�0�v�I@�ފА;��|�/fL�)�x��G$+j%.ܰNs�p�h���_3����Σ(�E�}:O�*UGA�d!���W���>��s�۔�Q�W��F�����^��\�z����Z�G������.�G��|�v�
 xWT�yL�&<x��,��sЌ��(�B�	�,}�q�:�,+}lF��p�-�-�O�	�^���
�w���W�6=B�f��7��^(��z�}�fp�5��U���������=�k7`A��'�����W&��;#Q�V�۽3����ڱ����+�}u([�P�����T8�A����^ַ������yЬ���8��c�O2�7���§/hL�Tc���p�i���S:��6g Ӧ����Ԓ
g㙐F#l��2�=�X����V�OIk'�K��,3ث���N��9=i��Y;�o3�p�B�c��Z����t�f눊�H�Ӟ� ���@6K� ��6ӉD��}U��o]}2��b��T�<�l�c`a�N�O�r检�-5�ְsL��(�K� �(ol�.Z;?m�%N�݅X-Jm8� c�L��T�m�
~6E%�Z���
�<�hs�W�"�w��e;�.Q#��- 	��xl1>p�]���.��m&�D�������>�p�;Ì���>hK����7S�Ťڃ��"XҚ0x������=�k�8c�o<m��Z�j�,p&}���EX�?Pʰ� ����y�ֻ�� �$�-}er��C�?X�� ��D}�h�����u�o�5�|aH˿�#25��1K�¡�~I��"�
����l���c[J�EN3��I8Ιw�:��_����f�@�*�-N�W&�R`<�A7T��W��xo�0sr��_�ZbbF�m��� �a4�[ރ�S�u#m��:,��x5���$pӢ��ˇ7���HSF�f>�8���s���:�Q�`㫙��Q��4��ҏM@sF��Z����h�֜(��(5v��SN���x&���wt��NT�&/���r��CYq
n���M��P���yц���^wݟP\��g�>_��e���Z���9+��e1S M!@�WNaUh�!�k�S�%+�&|4ӝQZH���q2SJJGh��;.Zk��f�oI����?�_΀�_- ���y���U�w�N�����:��эՏj�9��/�S�?��%�ɦ��5�9ERĪ8������j���d����ȯۂn@>�u�C�
J�17㾿]�9� ������������Ϙ�����U񩔟|w�1a�4�W/T���
Md�O��BQ�t��{3!?����H U���砝O>w1d���^�����1/�$@A)w�7s�Pex��B�vqo�l�����{X�(�[�Kz*(	c�T�h�;���G���g����R������T@��ѧ�U����>`Q71֨֙������i�nPEE��>�-)J�_z�C�(5gWW��T��t;��w��h9!�[fK9�xQ�Z��}=�sX���䟋7g��0���i�\�:K�_	x7�������D�b��eB�؜lO&���o)G$xUe��f*wÞ�1�}�ƾ1��Y!�,/Ĺ64{O�mb�|�R��X\Y��s�]�\��5��}�c��V1����~�����[��WbpH�Ư~{�!?��:����]��b��o���m�f�~��ݕ�/����}�A&p�5�d�