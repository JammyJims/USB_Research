XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"ܯ>��I�a���&�j���1��i�ѩb��(qx�|M��|O��>M%W"`k4d�W�ʹ%�^B)9�I{r 	օ�y\��̍k�	�I�M��q�Q��\���W��7�k�=I�;[(����@'^�ʗ�3�RC	�]�-(qWI�\������]z�)2l�#��Qg���>�v��MPb���ԏ�ю�����)��>���f�� ��Q����D|��.iO�����S���D0䯤�E>50��?����˃�0o<��U���y����d�#��'UbEI�`.���{ݙ�B|�A�2��/7��7�9D���2ɷ���ً�i
O��/�+v��eY�Q�) ������#H+g�k:U�Ƃ�[�I��)*|�4PHW����N.�O2rb�Vm l���Ȑ���/ɷA�(ll.^��� �9���N��c��[qɗ�t�Μlrv����DrL5qi�b��\��Ef��'a=�Ty�	�s�.�a�,N0�d��?S�7T��<~����gM�V�0�8�
X��cc���Y�]x��%�iǍ�K��Й�פ��O�ѳ�������C�I�
,���V-�g�suׄDφ*��Fa�I�cNw�8��֞�ةN_=Xzˍgevk �&?�(ֿe�$!ރ;Ӓ�����U�'��V*��m�p�r�o�ZQ����,�0��I�7�����u=[H{ ��1t��G��v���o������6�����#���)h�M)k�(=���zXlxVHYEB    4a83    1490�}�M<⮌~�i�(��{��v�Td�/��Ű_�O����q�Z�L�4�P��1��3�Z�.��ԀD�[��¾��z�\��ta1�F�í1O� ���% �-�9��އ�Q�gJ5���,RC_'7�s�@X5���|Z�06����������Tnb�x�%�NC��|"E�����+���/�0�͙Z{"���V�Q.�bj;@Ȫ��M��k�^非6Y��wg ����٨(���11���%n.&�
�qd#X]ya򔝜AA���z<�L2�tW^KfK����3>N�@3�F|��#�^0�x�EE*��h��O��.�/!�UD����!H���w+z���/����{ܰa9Xʃ�))w�'�p=`n����w��#��1��b���[iIeR�2����=]��D.�7#F�"i7v���30���7�q�:�MAx�!�a�,lf��5g���e��|g�G�����c��T�7Ӹ�(o�A�M�t1�B�(����)8��eH%�WgO�C��Z���f��>�����v%�� �(z�U��F�85?7�b�I���E�>>��$��s�شא ��^s�&��Ӿ�L.88���/c�o��V��|rR�2���B)*S(�?KÒk�8U�"@�<���I�U�*�~���l���Ia�jBQV�QS^�%Ư#���˓o^A�D��j�7\}/��Y���Uuq��)!D�i�Tpd5�Wvda�u+#c�w������C��Ȣ�q+��q�e��j�)_�����|��j�����O^6�y��~�u�}�����$cZȸ�r�;�ܵ;�O;�����j�}�GҝO�إ�i�>�`�3\�,�� �[BE���"�R��̃s�C��Z�!eq�rG�ܔ�g��쁻R��L�Q�*п;p�sbE���<�����)?o�3?`��0!@$����f����ȑ�;��9^I�.�V˜$�vvTW�`{�������Kp�J�+�e�^�<�4���"����-�Ms�1t��K�wO�$Qru�ѧ�fHP9�jc��a��)q�Q,�<��1�k�p��{��;9����&Ks�u�J�c|M���/�Qî��]�\����H��%m���C���Fk�1W!�E6�ʬ�Vc���|��^d]I����k��s�Z��0�Z��=K�.�2�Գ�� "���d��p���}$�~5��WgӺ�V3�B��AX���u�OR;R�"uS�,6��,NA�|��C"s:��(p"�ٿ���'�/O�dkDLZ���h��Z�{OLf!���� ��m�����E���G� �;JPT l����{c�1֊�}w���G7�i����+��,c���O�-Xg��)�X.�j/+�kZ���l�`_�q(slĴs�1�9��g�K�����&,ȇI˗��eY�)��N�9�̵��k�v���]�HkŴ���*�vV��^�eϲ�O�W+ ��`!W|sz�p>�[UY�{���Fir�"��܎~�d:�H�1O�C�v���s���*@�o�I��aC��!�
�Cc4a�r�
�|R�Yd���x`?�'������ܳx����0���S�>��sH�' ��k<��h��bw�!֏N��2Տ��H�LkrǬUJ�\�.��/��!�d�����Ꟑ��$��xx�W���!���\л_%�הm�T�"�����C����P��> �{3��/O�F�$H�}��$ ��W�޲h@N����H٠�Wf���U��I���H:[d����U���NWD��5|��*pc�^�{�}�m��� i� 7A�
[�}���Vېt�/2�;%���W��O����ʂ�IE�{�,ce�����Z��I)B�� ��F�+�۽���4ۧ�偾�{(tO��3p�|��#�q��$�j0�.U�V�z7�?�阆O���*�=�U(P�zL���cE���l
Y��m�
���[|}�3�)W4�勤
�%֓>�~U=���<��V�q�ə���Ӥ̔ݗ2�2���uԆ(x��[�1�O^�aNb$��}�Ӡ�׽��G,����C��S��]}��H[��	�Z����9�V�(�a�Ϳ���{�HYй���6_�T͚�zO�g����`|Z�֎��X�w�5㙰{#��W��#��y�	��>����$�<����=��YR%����Ybi��y����Wic����������D��AWB�mU�7��R�`�6�ܚ�G��!�K����:8����!|N`,zx�����Q-'d͍�j�.m7�A��6C���i.� K�1����9覓�qpS =ro�F�9C�H��4b�x��0�8���_����X���h��'_�~�U�˩i�`W#^	�0��Oc4��_�d�]��&���c���P�����w\m�)���>����"�l���{-iS{��z���#�����NQU?
mHp�F�?�k�-��c����(A���F����hN�'X$>l���q��:�4`��ԡ�]�WX'b����~�
�DF�z	�߀�v8lԲxںqz<�X	5@��a�k��X�]��1J~���NΙ�2��s��Ϫ(�^@k1��Q��f����,�L��X����@�����)k{!+	�]�w�%����O�Q(e�'�\CTT`�1��B�)��E(�a��wx$P�ߛ�%b#�jV4�8�'�p>�oE���u�mJ�_�QS`t&T��� 0��X��a�8�|Ø�8����˼C:ǅ%�#���1ƭ�xa]�Gc�.d h1	E���	 ��92�����`�-N�)7[�2�.�4�R��$���Y��&�	������=�Rƺ�""���Jsbђ?�8R�(M��~���қ@R"߃v����CF���$'�* ĳ�Ugc��\�u����О�X�K���St�ٜ��@۰�V�38���H�������էq2����q5��m�*4��ڣ\o�C��e@�Ϡ����g��8��<��� ��t���䋳s�{��v��r�AlM��ꙁ>l�9"<P�-mҨ���b9f��S ��,�����w�����WI}Bǩk�lFZ����E��� �=����?;υd��jڟ�2�$xQ
��E7�-�+�����B��N:�vF;OV>򟅊�AD�p�q��������L�X�������ŉWT^f:�����@����{[���J��	,�EP����C�Ĳ��C��6B�v������`�z�!��vyz�����2���߆@��� utR3! �:q7ЌM�g��{�u��Y�����g�&�CaPΗƲ��i'�U!Ȅi,&3�31 ��C�j�E]��6)B����&�?�߬M�vXύ��*WN�%�I*$e1#��,�E�T�Nρ3��[�*��c��>�ޗp�Ǽ4��+��У.���cl/2�j�E��C�����pձ�eZ�[@,r�/w�ۥ����*�5�x��[�B��FɄ�h=+[@����O�X"������ԇ���,E�<U��Z�q�|���s|^���?�Wa��?'�7�zȻ�.o�+`B
����D�iY\�z��:�]j�Y�u�c0�A7-�����s�w������n�������@=��N*��Q��y��� �.����2�������0���~�@p����"4�CA����M&͕��t�%���S9;M��TK�U��%p���3�^B0�Vͤ�i5/��:�w	7,Lw�B�����%�5ZPZ�|*�o\'����<�T%;7Tbr�`i�4��C␏����+��
�@oe���n]6�l��Uu]�'�1�F��o	/�N�e��עI�G��֎9�kW;�}CA��|E�biQ�G�d:�����B�Bu�A��v�����Ϊr�Csc�N+188��3u'F�%�s/���Vk�ɰ�N�λv���ߴ��x�{��z�:,�ć*�X������}N��}gM�zg�	�gE�_H,+<T�Z�S��fV�{��z�en۵��F�|5��.w
[�f"��b�vd�p{�;� V�;�N����6��.�]*/��������g��0���ʑΥ��]��֏�T2RTۀl��$j��ֵ0ޮ�d���1!I��ٶ��s���"�x�Xy�گ	KB�	�ʘ:���-i��U������{)#	�]X���6�Y'��G-�L���0x.��)ˉ�T���,"�)w�="�d���F�� *Ccw�;��"gҒdZD�Ԍ�-qVԑ�}��.#���gW��ЄH�K���͔� }Hق��}��ج�w�����T���s��\HR`T ��@/��,� ���3�T��$z��p��}D}�%��~L�d�ANx:�WMWT�Oc>]&�yi�RLA��.��b?���ݻ�JX=,3��ea����I��>I	���;,�E��s� ����J-�{d>��06��"+���`R��⻌����!Vȵ��K<#���=���4(��Ŀ3g�da�O铵���2$���]n�U���~�)~ʅW;1��yY���=?s�d��+�.�0�p4Z)!\��w>C�J���mȄ:�bz��DK�G�cLF˼?��vyG	 �AQ�ǾՋ𞰭��W$�wZ"�^N>�z��|�������&�4��@�!�]���a��/���ǧ�?����G�I�r2Ֆ*h���i������B��P� <c�]\���F��uA����֥�_��!�f}��L�N�m#G_c~���uN�ڶ�x�3np@}�������u����w�?��&���|��aj�����%��[^���9?[�d~��RF��x��֮MDk��9(��]�$����Bx�_�Q�v������Ų�t (�:[��hl�\5��Wv���L4VT���	W�Α�{RP�fhݡ����`��?@���5v�.o�nB챝7�#ם)�Y���j^
T�`�tX��l��W鞵9[�N��]����K����n�G�'�3�Jd;v^׍������N��5�h�p�/*vb�^.�;�����U�u�>�Xy5�
�S���x���% �#©�8Q��~��ڃڶy|RrN��|�bd$,�onL^���}�U��ռƍc�xN}�y�gUV���9Q?k�q�!W��vyG@�V�