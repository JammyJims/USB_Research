XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Qv����
y��E1�:���~[!k�f$d*ƨ��X�U�乊�)�]׹��H��-BC����\�6��9!T���u�%$�+�FT�_	Ɔ͐�:���e�a ��)�-Io�mR��A��3Tt2ڔ(BE��}��D��\l�)��x K�1~��\6R*¦H�G�_x+OG���&5Ƕ���g��D�uA��%���K ~��o�@�Lg���ֽf$2�x���Y����5� �� �jW [w���}f�-IG)��Œ���ZҖ�ۭ�L��l)�Z��%.4^7� g׸N�%����
�&����8��2�ԬT��B���4W;I�2��2Ŝ/r-���,yu�,|9�u����YQ~�\J������Z�*�z��3�[�]8k�m�/%�L�B����@.t��0�rW|�z�eU�Ȼ�-�r�������ވ1�n]0`��B�����	&�v
�7��4@�ǃ�Թkl��F�a�N�<j��IN����(I�[_�>s�r��'ѵ"�,@�ԕ�u�b��䍠�eQ��L�oa��ͪ�&�U���4��\�\�����F�ɜ@��a���ib��!��zt�c�In�_;6
&7\���E�߷o����)}z�(%�A�6��UŮC+�]�Q^>K�bb��. 1P�������Ah��^�B�֠���r�y���g�����hׯ�X�C�;^V%Q��'���Cr	j����bpZ0*�c��Y�"	=_~C���7����	XlxVHYEB    4151     ef0G���d;y���Oȧ�_�SLtX�^@�҂!s�oZ*��Uk%�D�v7��_��i8�/X �(!�\�I	EF������q*��"Z�S��z�2�	J�<w��\�ڜ�\���R���H���f�s|Vʐ�{Wn���Z���nf�v�m���6C�Pt%�y��弢��r�U�v:y|Q-SV���Z�(Ȱ�"!:�*t�}ix��)2��D^�M�r�x(M���^t[�2��d��KD^�k�;"Z0z��9`2nLW��a4�Yg>���p(lD�.�\����%���CzT.`�vb?�e��|�?k�ZS����O�c���ގ���.�Np���~�0��]X�;B�*��R^[Ⱦ0��;�qRK�x}`M�$8o��k�=��� �u��?�a�?�|��t�c��M�O��v.�A�GDC$�GǾ���?��n�-�	£�2T�'F(��+�ǝP����-4��2#H4d{�{0ZCY� �̓��t5���`؄���lԡ+�.��:vT����n�J\_�l�j��Wi� �c�|)��ޭ����Ѥ���>��Ek�k��������ⵛ>��h�{+��W��N-�N�`�:a��.=�.B�e��y)��?�km��Z�-�~�F��m���� z�d���f�ƣڛ���gu��
�zMה�=�3�<��Q�(�ݝ�Qy�/Y�7����T%��$V;�'�1X�9d��x�u��$�-�~.���ډ�S�g�Ÿny��u�􅳯M �x�W{�a�I'�8�r�2������$�%���P�e����_eox��"�I��dr���ݺV�OK�g���ui����*ȝ�����������}삩��F[W�*t��_^�8\��r")�7}nSP �ۥ&D N��ϋ8�����&���!���ډ6o{k/�⠤�[�Z�)�'�ݲ�׀���\B��Cʖ^?�D�dY���yW���`s�׆.$��p�.M1�	�A@�K42�Sߣ��kgw����BŐ\M��K�5�4%�jK�NՅ7yF����Y�z��f���`@�H��-;c~U<G6_÷YY/ڜ�T�II�⦭#0�g�}�|N���K�X[`�9�dMk��?~i7�a�Gu+��!\��FH���#�W��\��?vCD�N(�&���, ��?�8lR�t�f_9,Pi:��%�[�H���a[�o�tb�\Ð�KK��i�^r.Ƞ6)�����n���n����9a}	��š���I�0Ӥ�5�^��3��]8��g���`���:zܲ�M%jh��_�!�O(tS���U~C{��3�w�1���@��	%�h�_�F�/�^?
k�IY�cڝ���z��V�<CaȘ�I���<�p`g��BD,p�d�7�T��FF ��G�?���� 3�@,�q��}	���5@�m����$?ze���ѯ.JA�vz���ou�Mj� iO��;�$i欞�������
�RD�s߲'7/��Q�k,p�A"�j�5��	���Ʒ,��2I�B���H��T�_c�J7$�$%�9��G9�^1kd2m�@S/㑿�*���-s�/ևi�@�u_�=�ȢNQH�ߟ����B��v�È�]N�WnqX�l���w���j{�����*�b,:����x��gV#r��i�k؂��C��_�=�H!�&ά�OCLح�K�o� Ua#��_��W�Q�W�37��F�B���2�������g
(�z|Ăi�sPw��m�]�R���/�
��j�d�1 � -,7�q��]�?Z�~�v2�{�Pf�9��|�hG���L���Z:'�����V�)܂��dHzSN�\�	�0�U�L�y-�o��� ��l�O���-�.]b��[U��}j��V��"�ix����]�\�����gkT��G�����!n1%�s?L�w����@�K7�w֋/ﳜ#d��/^
V2�V́]�8��~����K@�u�9�jY[�����VF\&�E�"׆���c嶜� 1�FMS}A��@)�d���KԢ�m-��ʷ��I�	cX���d�$�GW,b8:��2����^�����^�GS���?[8��s@�|q����_'�?�ޑh_���j�L��u��E3r�ī��������ў��*+K|e�T�H� ��6�{��֏)��V^�Ia�z�[�v�2i���YiWW�~-���qϠ��n�6��xo �dj����5�O������ܧ_r�`]t�X�F_lrt\Ff��߹������>Q�a 
�Q�tF�3ԗo��"���ukh�ty�'�"����cC�5q�IF� ���_�bt���^��(����?�$n���Rv�^��j<��X�W/#j�����â��Ђ�!��� ��4�d*,=0ʴ�:���ci�_��
�4�ȶ���@�2��")�	�(����$ʇE˽�aۇ�rʛؼ���D�)�����!=V�⁒Y+��d�lqŸ���7˫���5@|l�U�^WS�M�)�;0�n%X����w�Ѵ��Q��;(bz��к��zk�G��]���1��\� � �ջ]7w����w�~K���5B�>ES�E( �B<q}"P�Lk��ic��� B�V0��Т=q�t����e$�5�LC��m�h����O�-)��C2 �A
�����}�k�˖H���ĵ(��6ͯj��n�N�N���Z�w&�'��9�Nɏ1�zmY�7��	��#3�b=2�T@z��9�r�W���fa���Uo"� $�[�|��ޖҾL�gi�ٙV�,ǐ��g.��m�P��0i&5�o���*����X8�e'h�Ő�n�X`C)�:�U�	����i'�_�e��@����L=s܂�ԇ��QV�,>қ;"Q�5�À)��.&~�S4��EF}�f���bmی��O�����d�>���ff���bi��q�n�%�)�ʩ#��}4���}�i�f�b�5�а+kP�;�"�wm���^��+=���\8o�64Pu�p�o'_M ;=Eݭ,[���^�>I4��v�C��Tn�����-1��<K�����-+�{[����}^��W���#�����p���y�g�6Nbz��Y��bvbbZR���ŀ,�库�����'q�/�.��_bdչ���ڶӶĀ,��}mچ�ٸ�z�ih��
�A5�E.f�	���)R���.�O����p�,({%�%'9��O��Q�.��<�}A�O�tU�#$��3�a(��â�e�$o#T()�[v�ZY���P�hѓE=��$3���gn_^Qp��V����f�^Jki�Kۚ���]���F%�\&�w�����&Y�o�8�X���K���ƤUL��(���e~��KK����s���N+�W!V7�� ڛ*�^��?soMe�#�l�w}lV4x�DُJ�P�)\1��iň�*�%�q�$��(�,ZM��H ���-�U�J���T�BG4N9��[ !��oYL���v��<f����JT�*�4(&4�N��:�D�Sv{�*�)h	�T����Y��GP�-E���HQ���=��`jD%�&p7��g�[����@�^N�Z8��a����ߋlεЧ�ގ�zK#�>�j��h�j�!X�c���=��RH�>�Ӑ ���T��ot2���I4�c���d���?V��m��x)-��\I��|-���jh_��aoF�0�<���U�YUS19k�n��i�?��������Ղ��JN���#���r�*��l&�s��d������^��?