XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����]Kn`��Ǫ�I "tO�n���D&�J7����'"�b.��%�LHH0P	�5�\O�8�X�5X� �~ V�c��#nwϲ�R`Ʃx���L[Rg���;��c���*0Z�v�|l:ɇi�#_�U��֝��R�:![���������ϳ|R�-�[1�i�BWR7&�������j5���W�#Rb{s`@ɷ���;��m�e`<}E`���}�v��X���8�zm����*h&�e��D�j_��%l+��>�+D���N�j����v������~_m�3����ԁ��yY���2J����zB��"�#�X�(���O%�$����1õ��O�Z������Ք�u,rCWK �U��
g�AB�0bwq�Жn��*�7W�d���+�C_��<��*(AS`���I�U��?]S�2`����6�"԰�tyru��p5��!�A���y����	�:�k��gx���e��I��YV�=�9�>�*�a�<y�x�E�/��8��,��5�>n� dB)��%�"��$\ao���їm���V���E�R����	
��,)_�5G-�����AȺ�?��-sR
	����j�wvq�n����L]eA�-1:�^L.i�_-
�q��Pǳ�}�)��<����;X&��)r�|��gP���*����"OyV�L���l)���e�UMT�*?���_�S���[f���ϑ i�1�H"�l�k�P9<7fHw��P7�ВB^�6W�XlxVHYEB    5bdb    1960��Ġ*��0�/(s]Z�����bmE�)�\aB�����x����xgx�3�>��EP�F���ڢ�,F�}��
�"�ow��]�-��ѥ�*^j�B��0�YZ־�AY@|��e��ӑ$�_�B���qt˶��U��u$�`���~�~<~��k�iƬ���A!��cl0��2�cFAX��4��0�օ�?ߩ��^�["j۹B�ֆ��,RE�B�̈�%��]�[��CR-����+HY��0�U�?�D�C��ym3�:��^F�<L>ݷ���M�Y����,��i:��e���֪��F��y�;���ho��-f���JS|ۣ9�����З	-:�Zi8��V��k�F�^�ΟGx�:�g���(����	� ��j���>��#�xl¡��h�pu*BV-&��E��~BjH�q�,�)�n>�S�ϫ�C�ƌ!��YG���9�f�o�o||#��W�w����b]%oHR�buU���&�#}Dr!W��F3���#���*�'��DGWC�Q�
��g���2��U����<��M�mnna��p�#%��Ps�߄��}h�D��[78~�~T��u��{��Tl-�T��z���+��F3>P}���vg�?��UYb@��hL�$B�J9��T��X��f
)�7���p��h�*	˹��t�A�d<�U6 �ʭ���i#^q�ٯ�I��������-�O��Dp�8_?(q,��v{�sH`|W�(��i*�i"�C��BH����b���}����
rܘ�
 �Dȅ�t�kD`��-�+�X�-�����d�Ô�9����֚Kݩ�>�<�g��Y�U�Qţ������_�L ��L&P':C5^M`\���Ŕt �hJ�=�p]ƲqA%��y��K�U[}j%D{������,�o��:ED�Fw?ꔭ�i��l=>V��7w����˶�-�",@������l���
�*]�߽��r���} �H�9@���spݛ���[B锏@4ϩ��__k"�������b��,�z��<�&�~��|�L�����N� J�[5K�GMx��AU��B�!	�B�a�O76#�v�j��~4k�Շp9���F_ɋt��=1�FLm6�nI]�x���1SÂ��K0d���XrҏU���F��/_���e:��)
�֫h����';��eGQ�@p\G+A=��ݐ��}M��g"�������ɼ0)Y!S��RK�Y��_��`��.w�g��U�J��	�� Ә��[�1,�'��HrL��0���]EB�8�*I�G�ahil�����}
�D��	{����=_�sU;_���h4����8S�:đG�6@xyJf7lc��Z���bں�㛾�9�`mμf�F�0t�F��^eh$'��� �/���)�X�}|�s��vQ1R����T�NWq��}1Fn�H]*s�^�G��(Pޓi]���D��-��ht߾Bo���Nm����~�N-�F��E�?��kM5��u�"~Z0�t�\��Y� �ʖ�]D��,���s�#�z�]$����j� &���Y�����R9A�ZUF�釆Ϧ]��L�����h?:����ZVK+�w,?������C\�U��Hɹ�͔Εq���u*\�	���0[b�H�s@�Y��N��g��?�2��F� �(g�l��=i�64������B�8F��W�ȧ�i�'���K���a�V�(�o�}(�Y����r��/�ܠl���S�s�-�/XN�'ꅨ��[���ҳ�:�傿�Z[-�~���n����y���(�^c�,\�����1��-��w��\&�z�h�b@�� F[g֐@�Ĳ�RR����XW���0�,��R����?ؘ�[�F�^z�$�R�Pi�ؾX!x�����fζ��z'�$�z�if��Â,�`'��\�m��Y��gHu�G�":��GQQ�����Yr�9�F��!a�OSU̓2
R�J	q��ʼ�Tr�r�E�xq�w9A`��E�a���eƏa�8��J	zB-;�� ��N�~6���8rŐ*�O�G\�D��S]�"�Lg�/\��Y�,%��!S�_��ꤡ�e�U��O�S�x�hφ����BI���.����7y	�����TT��_v�i{�Y*�B����bR�!�G�;T�
�����@����$P�����}ȖG}S�ۼ�a҇�6ʌ:߬橘E)#�i/���c*�*�+�[��i��A6��.���!�W�E]bq�ײ�����U���<�'���k�� �5��zy8ǩ�����O�MW��4��en ���e/J��X�'R�چ�E�$D��X�P����õ�ļ*�p�^h�rrg��h�{=wS���l��,�e����E����i���4���?�ƒ�n��;�+�<��8�B�mN���V̓9����<����@�3�7�V[ I���(�Ch��8�� �+�BŅD`$� ���;=7VĹ��X
��S��r�h�R�lYH���M�,�%���-i�GJ�j�*�qd�n��<.R+��#JOd4�F��m1������8My�BZZ�Y��SȘQ%55LI�Z�^];4K���e�}��34�V���@Y��E*l�1��^���5W0�~�����H�s��f�%I�����RkE��@�J��2m$Q�7���K����m��]y#�+��򩞆�=���k}�VH�]`���F'�w�쑍"��q�e.�h���9���?�1��1tD6�ӑ�-��J�0J6?�v�J�U�7�C�TV�k;��<�I`�o�[!%2��E�ND��BG�q�(�Oj��>G��}��� �@���\gxVMQ���p�����V�T���\3��=͈Z֝[�V+�!��4�]!(C��
�V�@�IwЅ3l�K�yN���؛:1�'��Rcgy��{�w�e�4����dA��Yr㳈�E�b3\o_bmш��U�l��m�hu�Cj��%y�64O��1 ��A���Zຂc��:b:�e���%��O�uU��j:���o ��_U��V�Q3
`����1��.N�4}Ws-]�����4ϨD)��o���_��Q�<Yg�(�>�h��p�I����Ʊ%9�Z��H��_���~Hiwiy�)"[h�ҝ�����,os�]$N�S.��Zm��kC��@�o��á%�� ��T8k2lA&��aY
��&_' A�E�r��3���<��1o�p�����Z����i�H��$\JM�`	¼
�� �[�4~���?d7;��ϡ�d�»S�����W��8���*HL�J?���5�."H�TUh��#�U��f�mtq���ZHU� ��J�NU$��V=e��*C�K�,����]6Y\§d���'h(%�f�r�9�L�V�1ԩ: �˩b��B��yF�h�dA)�U�j�G.xjvZ@��K�N檎L&K1Hy���K��-��U�|�aM�4���;�6z�/�z+�,�N[oX��f�ϖF9�r�Jzq��£�7�����L]��	聟Oo��$W�1�L3���0G�C�VT��M��A� ����)p���CT�b���r�w򆤝^��~�E��i�LԔ��r��m�]6~��*7��4�e���M�����-�m>�L���KlZ��Nh���&0\��`�+f�\ǲp��8
�B_��h����hS2*5�)�:�R�ˉ�;�t���/w��[�m�w�J��C�{�����8l�5���cj�&:��0�e��C��|�m8���3�b[�S��_�/��	���R���~�HB0��>ӕV-�ѯq��|c��Y3H|ۗ��%_�~��u|�\���g{�=��ޒ\v~�-�����(l�C�T�@g��)3o�Lr��+��I� �]�#V�����g���յx�۩!-;�$/�(�*X�w�r��E� ��<��$$m�!�>�A�p�bCNCBݡ��]̄a/B����lS��{-���}����'�>�7�H��.�z{fzؓ����#�+�r����O�`��!s3Pa� :S���<E����b�������q�������`�IC}
+"���m� ��o^kv(׵[J���L$��%\��=u�.$�z�W����W���V؈2.��wW*c<���l~b%ޱ(���ĸ���R�
���M�|�R���F��F~�]"��7A4��3ܧ���t�<zfG�ԡ��k@�����X�2�X��W�I�6&q��>7�.���D7��4�nEE�C2\��� l���N��b��QZ���.�j�ڰ5�v@��mjp��^����A�$�L'�,�L�>��p�o��_
�},���MH[\r�ڎh?`��̗�� <i�]J�u���"W���ɲ��'>W/HH�@2w��Ք�t2���nY�eJ��y-E�Tn��,�[��Чa5�[wU9a-���mu����=*0U��Hb�'6v
͔v |5!��*�Ū) ��6�^={:Y�q����W���H��!c�L�'w'5G�Sڰ
oh�l��H3�<y?�PV����h��u���)�&m�CN%��L�U�vb��dE*���u<QZH<�o�P�n��tD,vLze���^���LX�� ܏��/�L�K��m�_쀘��ZV~��~l�����^�򎲠���d����Z��Q~�*�
��@����G^�A�	�#�4wHqF�<㏾�߶����_k�~Q'��+�d�	Vm���қ�J��6'���a{�`{�O�ЭF^��`��صIA ��g���驇Vܹ@�D�	�=�� �иG�{Ot�z�,[�eR����O�����
˭[!Q��]W��Z~��>���i�'y�|ac`'��nƗ�����7�8d��H���2^�wX�&mge���JP�n�	X7x?!ND�9�Oo�B3���7Z�ϝ������?@f�6�!t:�����ﾉaX��Xl����eW��k.���hN1y5	��s*� iȥ�"wG�P�@�HK��}rE�f~���Ă96]S��z��6	D�Q��7�6=�R�dN�$�xngF0�?�ko��U��7)!�r�nR�K���AIcr��ӍT���%��n�jr���o$8xG{���&!a���:����Չ�&��(�]�]��� )*Ex8:�7u�T�uV�.G�W����v����������wV�sE�Nϱl |�Э�Rp��|B+h�,J��ㇿ�
��:��U�R1s�ʷ��N�>��n'xu����ZV��?�OO@�{�V�9�K�\�'�%��$��%N�� �@V��o�]��x�b�2&笱c��w@%�a���Z2�6���
����#� �%�ot+�m0�*z���I�K3�g�� CbH�ս|\�v㮳�f�󯁂�&�����v�1�[VI�܌h:j��wY3'���M6����tb�<6�7[j��QM7r1����հ�Q���2 o`U�暮����=oD�-e��Dƪ຋1�t��'>u\�4��w�$�Ury'#(i��(����-~�|"�Gʫ�'�]���֒]�����l�~��$PX+nZ�b��t�j?�a;�`/9�Le�dH�+*��1�֐�F(}�~%��Qs6���e}׍&��i�z���P-'a'�Dޟ�\{.��Bh��Z aM���������q�����K���zqm�j�吏M!�+w/�0��/{���$�isNKN��p���>�N�@[�+�O����Dix�Rq��쪬!f����,t"�^I�Ǳ)����ef�
,Ϋ�)�^39�A
}��~���weA�V�7�F`mi̚����M35�&dCx�$U⧫6^ �%��g{����4'�R�b}� �D������O뗗Þ[vqƙX X����!_4�*��1�J��a��B����lr�{/��/�V�$*����l��ί�#���j33��2]*��B9 �{C�Rs�p�{�����Ms���+�ި��=�9�cFI
¦� -�AO�T(��aԦ6��[��:a-D���:\���z"9sCE��;�<��GlQ2eע|>�1�r�"���H�k����4�B/�ݫ8e�k�2�d$c�jg�\���j�x ���R"x�DA����-�G?��?���C����۲�r/h/�(�G���2�V�.9^U���V�-X�+��~����~(,���5��2"�3'����c�C`�rE���G�+u鰒�[[�|�8/E@P�6z���o�2]�x�!�{���#؎�/$Fӄ��;�H��!i���H�>��rOx>��o����g�S��@��U4�Hk�ab�p�Խ�%�ss5�U���2ȭg=���ևB��x������i��cq��8��0\��QR