XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g+n@I�<Ba��}��������g������j3;�۔���ET�)L_�|+�3�B��\�mF� me��d���-!L�~�oR�F�Hc��Ż�g���5�3*�{�f1E4��!,��-IJ@WUq.�q4�q@p�'�(2ӽ�NNN�Ĩ	V��T�0S-(A0��0���I0��(F6��Cp?�[��	�8�}�����n]*���b�������i6`�|�=��[+� wVk-߶W��31���dY�|��kd:���]�tR�;i���|;����aĨޮ��ScG���h��8�'�3�e1*�hΕ������� ��m q"��πSZ�sP�+w�eW��U�qo�q�*3cUx-z�[*��Xi��`$H!sBs�Œ�^n��vV>�`������@u��Ye��ϗ�@�M�꺲u�K����<��g 3@�hy�A�s	�1��zI0�t��i<����k �H��N�����%\��Y��3�*�he��eLd�L%��7Q�
���C�=����\;�m����K�U�Q)�s���q��ɇ���6�~Ԝp��yJ^B�?�;�����L��#���Z��!�xiU�A��m�+'0�M�������9�_ݤ��C��a���B8�7�������d��x�$�:ґe�O��h��>�6c��
���6F0��Y��A���Rpc�z��\��}�5�� ��]^�N��>���%�ᰑgv8Y����T���L������o0�\yq { K[�!XlxVHYEB    2ecf     d10$�rr�n��8m�xU�U�/4`nN�;� K联�:�q�{������G�$��ӯ��,w;��@tL���D��9�A�b֎_��L��ɮݸ�#�*^kHÂ��\��4�{��̆���������_Ϯ�L��Ku��ެX��=ߺ�]�m�$���B�B}r������}�߮���{qߛ�1t
27i�m��s|[���1��Ɉ�Fxs%Ȱ���˳Ռ^��9:�ق/�~��C"���!���z�_�C@�as�X��R�S��ֽ����u���1�
��|F���Yvk�)el��9�D��1�QW��O
 �f�#X,��l��K1f�ڍ�� /4�_1�h/d��,(L|�J��ܬMZJ9��v�l�Hg�$�F�W��H�/�Gf��^��zf���4S��`�K-K��猉�ڇ�7� �~�@w�ٮ2��>W�?k�hr�-��ܥ�W�QJ~L��A�gL�8"xd�5Հ��\��~�u��Q+n�k�6'�É�k�H�E��k|˾�M
䥕�k�w�ڌ�Kz`G�SA?*	5��&|�E]�\x�m6%΀��Pdޑ$3Z�?!F$w��-���KÞg�;��ڄ�������V��_Ox�f�k
��A�qH>Zؑ�`�s��rg���Q���/E��ܧFu�5pΕ_���;[�Ӱ����������O�P���)���ٟ�ڹ�B�S]j^B�etǐy%^5>eC�����Dˉ(~����p��H1ĕv!A�c�1o����+��ڤ|��AAv=�ϳ�hj>$��,Z��o�W�i�S&MjT��$�	�ڀ�T�Yߞ���2$�C*_���!�~Uܪw��<�j��PAҶ^� �@.^ď�V�X+���n��>VdݲOLDI��.qQ���޺�)���./Að�Ofq4���|�[f�)мPCA�6u�Ӗ�";h
���yP-�	������_c�?��S��݂��J�Yu� �?yT�7Ul�O1�F����0�2/"��rψ�$�8,�%���%��O�[h?���i��]ӕ�j:��QF�sf�!����Lo���G"�����3Q�!VJ�H�1`P �۲�R<Y��]r�G/�t' 	qfSr��3�ve���#>J��]���r�������D��i�����q<��B>�)@�m!����Ԛ�,#��,����5��x����bg�U�&�핺٤����1Z��u;Fx�{���?���a3c�_g�T��2��{�{�Ԅ�뭒�&��<z����Ds�L��`���M�ƱJ���/�H�� J���-��Ɩ��� �j�����C���C���;m{H����v`��F=l)3w%#��)��B�}�l���b��d�!W�G<gDG�Nb �
K{�@̼dz����MZD��*rB\��~ ���_Um������s>��,T��=��*�r��oë8�D�T)Ko�&�5W|hqD��9�A�&�(�a3,[l���3�hS��ۯ�9ePeG�0NN�h�R�����NI'������O��zx��@�����'����5�������6$��@1�g�@���p�p�9�!��7����+�^;�v��,w{�r�Xz��}�g�W"_�Q��� "�r>g��Ьr��*Wr��/��V���O�iS~_�?y�� �!hWh;���'����`��
�,���ŵ&�V���ْ)�i���m�q�ȫKz.!��*_�����#��p��}�T�)뷠���Z�xC����1�3�x�$w�vB����P�j�^p.������E㱓]N$B�C�1� �j�	��/k ��q܏����B �#CDzCN���71%֪��~`k��b���8�l85lB��VxG�s���@�9L��{������;�Y%��wұ�릜>��#�3��X�܅���܂��g�a#�2��4�iyX{�j�@j�Θ�?���j:�� ~m��R�B ��[:��P�&����=S�?aa�G��z�̢��\�:�I5�T�}3�'��,�I���T�)��Q��"|y(� ��hi�v�_,FH&@?ClA����o��G����?�<�_�1�����tU����a�)��4�!9����\j���=ŭO���`&�:�������"s1z����N�q]�W{-�8���t��L��eN�Ҁ{��H+�Uj]� iYp�H~M�\�O/;d)�N{|��)˶W7�3���a���M��Do/�2�.r��%�V����J���P|uX���eQ��XӲ<Rt�r:��I���0`�1��7Q�t�8P�伥�L#Rt/�$C	�f�dQ��c�2��f�i���'��E�d}ތE{7�=FBY�>h�i�R,1�,��g$CaZ/�Dx��/�)��y���z��b�ix3,pG�k'#ẃ�֮@;5�9�����&�u��U�J���1��ĸ�"��t�FU��(z$"4$�GϏ�/���ԛ�-a������ͺ��kx$�}W��mhS�H*�1��
�5X��J���� ����峤čQ$�i�'�c���;�ì�e�a�,��x6�[ 
f�P�b�;I�tᚡ�ŉC��G��6"˷D�Z�0`���������7��L�j�*:�ߖ�$Λ���Z@���e �K������|)�Ɏ��h��[�5UD��l��ca����	���D��MB��ǔf�[�&���vP�E��
"�A��Q�&�φ*'�v��0�Q,��i�P �P�0���8�9��y̒�������k�P�^�+4i(��'�,�(�	q�g�*ThJ2�PƏ�?*��e�g �����>�-��R7�ϥ�U8���)|%tu���H�J;J�O���_��
�j�y�(�(
T��M�Ѵh$.�Z|�^P79�����'�� �X����ZA��g݈���T5
i̋.�MJ4�+f+0��>j�������=7�Al�k�͇��R��$�oS��V[��LF������Z��vn������&����i�f���|ߖ@��o��
�Q/��v.�"rIɦ�)u�4�a���x�Z���X�P�i�V�I���Ҝ�]�>�<�0Xe�����?�f��@ ,{�v:V�z!<[*䶀�H��C��d,o���+�w
3\�G����ea��3�#��!�Q9�m�<a'Dc\�ؗ
7���KI6��ڻ��~l��ԛ���=Of̐�ЁD�����Fle���.�AN�S��!`û�9~�2�8�%:��ԔD�����t��T7�`@
��