XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S��Q�B�qz^�p�܂	�H L�Ȓ�5���V��δ�	�9�[���?����u����ӭ*�H��cϓ��R65H�h�������@���hz/F;����/"zl��R�Q��K�z�
Wj��4������_�	���N�x3�a|�]#IM�=Wz��b/tu��-����d]�,%�8/�[ �ς�3�9L�ʇ�Jf�o�s0Cu�`*M�Ih_7�9�W�d�,O}aO�h��?���T�W�٥V�P�@��Iб�B'�U�u~]�}Es`�T�}ƕ��I��0�e����<*bW��E��H{� �K��+P��.tI��w��
�8�����e�?;P�< ޭ]=���0Փcӓe�
�B��D�J��
�t	 d����?�����7��a�^#��������A���A�!i�6[�f��W�'��U��]���Y+�����0ç]o�(<A��L�S�ꩉއ�鏌p2�9N%_��Q��q�jΤ���̼ĕL��4 ަ�AA�f�I>�7�w�n�e�6�$�~R�z���!'���=��~����D��J�-Ǻ	�!cT��(����[��y�r�I)�J(M�)^�ֿh�N�%��MR�N9$�E�c��I��Ծ���X���w���Zµ�Xo&̆��w}@��e�	�F[�2�W�樆0�\-�uQ��u��y5{Mo�e�J��'���{ �e�Fd<� ���8�|Lw�ZTJ<���Ycy��ֲ��o_�@r��XlxVHYEB    3a42     d60)c��pvϒZ�C��qm���5���p'뗎M��O��A�؈9���^�Ẍ́$�(1�c�a�o�
B["���
ܬO_|kG}`m�R#بF�o�J�\�k<J��ę�Q�w��E~GKz��a0,?�ȐVO�Us}1+����G	D�<ɡ>���ȝ�٧��2�L'bd����U¼ ��_�=�F���k�@FtFhL�M�%1�E�o�Ѽu#��OD�$.|�U���l�35��l�4J�p��2��k7�ɶ4��B�vaѸ.*'�V����nK݊c��<��=�����8�0��K�.\:fi�叽d|���h���{�W��f�A����D�����P�V~ �cɂ]�XC��RK@�W6�s"��(�e�n�꜄�,vkb9�'�u�����,�v���S���Z&6���|N��K���!Ռ�<�K�����Bi_(=��.���bil�XygI��w�T\�Q6݌�5��j�)x�s�[��oC�*C����	�Zț��$џ������s��T���E{ÿy����R�(��]/�+�������y�-�>���5�����3D�0���-R�i�!5g
O�����J���E�C����kH�m�Jg���&�������:�%��Gh�[�s�_L�6s���~ ���t���ǹRxd�m�&��n�X�%�L�n������av�$����S��bF���_��˾� JZ���`w���'oa����S�W�e�em*q��	6&G�������y����Ⱦ�g�7��¡�)���RQ=~��u>hMu�c�#���t^��x̂�|����V��21Wö�I1yt[lE7��:E�'�d�럼�<�&F�s�(�(��a�1�����W�����r�Ѳn��������vA��WŹF��L�̣?a��J�(��2���-���,'�Qٛp8� dUP�nva܀՘ۡ��%�x��vl�!�[84r��
 �c2��r$z	�p:��y�X9x�ji��D[�I9V6V�S-�o����r�����k�]�}TCe���y�@{2�xkdrP"��b�r�_e� `[��(�>�PM�,k����k�~ڕ��r�P����F���c'����}�;��I����]n��[$���e��ܩ$_��H댴� Й�|ښ)��ӎ�\�Z-2��t�Ľ��e6�]��x
ݚ�oHNm@<������Ć'�/\�����r���3Z�(�%<س��	 /���/���hH��T_�V�:�++�ٽ��?�W�>k��b}[�my�)���,���p�����X��(�\~Ò��D���R���}�M���
]n���q����ErR�M�P���Vq[P�Z��,e��w���l��=<;Ndy��2��5ʯ�\��IX�t1<�dr|2���/�1t�����W������#�� mw�2�)��.�B��q	~�J�O��=@5h�`�A�o]�и��а���A���OA�va�����wm�(՟���5����U��y�6�	+�����Z�g����,c�]����S���I�L��j�|RM-��F�c�
�.��N��	��:/D��,��68e,���S����c#���02.�9]�� V;{сR��!�`�5�͒	f����]a����y��������Zs<	���� f�=��W8����'0�s�^�,�r��ɰ��1�T���3]:@4��U��H���1��nk�7��9J@*��~!���W���g#�I'��R�LO�ڡ5]Q]w�B�
ۼ�$���-~�4Z��uuۑX
ZlWS�݄|q՟��h���O�Ra+�\�}t7
�N�<!�����t4�퇕�DK�������T�:�Q�fz|�0����M�[�w8�)�	]�(5�R�B��phg`BI~��gܳ�yJ��-&�[߿\,�hW5]���������4�1Ν6�C��I�ı#�}�,������ֹ���^T������W��z�N:[I�tpiW�jB�e!�������zK�z������@�:AI$U[�I)��:@&F�Ps����I�a���]���`�~Y���S�x����d�؂ܟ���)G�|����߁ǿ�9SP���s�l50����Au�H䎠�,n�p׹����� ���"'�f��Gl!Z�K��d���R$a�Vǉ^�����8���i1=Oɿ�yh�����:*�pO�1�
�R��Wcׇ�~S�Brd��m�3I:!�)h�#�w��q�5xC���V�(R�+k�]̲���̟�L�36��#, >-��=-��~C�]�ҕf�T�R��Z�X|e�7 #�������`�r�����L�xVm�Pb=X�du,�Mw�Be��߆����)ϓc� Avp��9��<�}�H�>a���Q����>p�%�Q��W�)t����/�j�5�uV��\�88�ӟlF���}:"�YUT����p��ۈJ�3ǳ�81����d��nG�Fv����2E���&��&k/��QK����Rn��q�^Ô�1�6qQ%��(-�Q�Hp36��~�y��ߖ��x�Sڈ�r)խy����}@�L�L:��7ӯ<��jl�K�s
y�t��d�?_o�S!8��ed���Bh�$����s�
��3ˁ��i^˔_����$E�#�d�i�k�$a���"Q���M���.�ߥ�QH�x ��!��u���r��3��q*wI5��Ն���e��Kq�=�Ha��M,9]�e�&7�C��@�Y�� n;`>9��tO灗0���;���SÜ6�]�ь�o���N7uA=
%@� �a����r��w=������N�$�~yv,�<sU1�����������V^q�d=�HL0{���<�Uc���y����$C����S	s�)3�b>?�C&!������bT�	�&{V�@"�|�1��K��q1rdrx*ڟT�ĔbNu�����kh(��7f�6u���d<�vJj7�Q*ຌ����<朲ZPn^����V"�dN�Ȣ�9=w�y��Ą��|ٸ�q��Ǻ��HB'�Xz��|�;�k����ڗ=iN�����Y)����>ȝ���BYo����,&����~��T�0�������{D�X`�y@�5'JB��8��8iuN�VOw��gh�&|M�*�o�G�b �YdeNk��c��f)��f;�V㔫^�<����b��yBwf=f��<
���$l��z/0Љ�^�Zj.���l^?���¥�6'���a�J@XG=96q��{����h��d�B��ee8"�Ȟ��Wǡ|p�%F%�=_ .5��J-���/��hX#��Ϊ��IV���^8E8