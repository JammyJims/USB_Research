XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_>��@��C��͖t�Ќ�p��n��AIU//����Z1)�.w��V�)�_kT�����յ훰�"O�hڳ���}��b�M#�رM�C:'�Z�r/�X�h'���}0�f����B �����[�h�SA:��D˷}*�4h�/�+� �71��%�ҼQg�y�7�c�ȍ�9e�r���ڡ?���
���5�Ukv�
]|)$dĽ^����.N��,�Ǖ���zEF�a��f��/�39�I��tஆ����a��ĕ�w����]��}�h�M?mR�E�xj{�0��݊�g��5{>����-��^��|n35O������L�i�����K���{@�JE3R�����T�/�8���O���*�<ߣf�V���9��PqN�ʔ��Ή���}��J�x:�[qL���KMcI�A�{��>���/�n�u
���s1�Ʒo���k�7
��,���`Nޓ��f ����އ���O��N�쁕i�0g���Q��q/ӗ�g=	�g����г���}
p%=F�ft%n!"��N�Z?uwp榻DWy"����tR���ۮ���q�����Yp/'M��\����ȹP�%� �m���W�J�,G�"��YP?�p4]Y�>���MNþ�]T{=&�u�5_z��HX��%�������I�j�{^@�A�&�-�F'��f}y�x��ᖜ�C���_u��f;���I��+ߍ`��������<���n��2�-?��S����1XlxVHYEB    238c     bd0�ʄr�#�c� k�=1xϔ4��8n�/����cRK���F�e�G�U�k�p](����r'Hp���X{!ϿT-�NM��࠸[���g��F�JT �Đ!�����Y�öe�ޚ���;�3���q\Zw�1k�Gh�y#k�'��Hϲb&!$��k��Tx��65���(�n�Փp1r�7T�n��F-hl�P($�>+�U��H�ŤX�����.�D���m�ZK_�2O�D��)���פ���q�O`�	.�]�<��)����O���v�<kt Aa)fIkͩ.�ŵyaŠ�<��=�H� �獩�Gyz���������{n�o���j�
o�AZ3u0��}˾�C��n�l9vE){/��x�GX��t�;�"�=lq�wч�i��߶��|��íN���ߞ�����_�λ��ב➴���qG�P��*c}/��^u�|�wz=�,����� Wl�f}���JJB����J�:1�?�����%QǱkQ%����ÌʋkRu�;Di�_u@P�����r
Go���q��IxP��əDٸ�o�,F���B/�F]����ǽ�=��o��O�Z=b'�y�'JX޹���!`�$�)���Xvٲif��~�q��6VV]=\k�@I˹[���$x���$N��m`��1�q�*�ӥ��ڍ��~���|���)i)��F#?T���p��K+WD;�I�2��t��/�a�˪P����R.�T����F{(���5�';7�gz��]��v��rJ�N��`0��(������.�L���]�η�ĝ��F<Dt8�ez�y-
�� ��UMK]���^��]~��i�K�V�����l9R���b HM��1��(v�9R�$Ybۛ��� �m�\ ߕ9��-Ǭ���-��]������;���՞�7mDBD�y����r�^��U�T�#���s�Ps����-x$��ĿP �c�J%3������c�1���*a�B��B"�����g<�ۗC�T�N�"��i��_��GZ0O[7_��F�)W����V�y���rqߍ�vd� ��� 7����2����w�8�����]l��j�Q���&*wNu5�E�ӵ��
1���܌@H�0h>^b��� T{�v�(��x�K�2���=
�բ���i�%k����p��XZ����FE&�T�ب(!����@G%d�#�V�đ̜��Oǆ��̿,3f��л���5��P�s�"�N{r��<����MA��^r���ǰКT�U�����T�����`�Bx6���@!v�Vý�=p��]$��Z��~3��(��H?�;�����W��{���7����^b0��{p��-"���O�hY���E8d��Q��[x_�MQ�xҴw�Ÿ�&O��H���g?Õ^��U�C	�HW�un`�!�D�#ަu��I�zI��sy8m.�nʻ���䉐��\]r�x`�'���N�&St�Л���n��Ӓ����4;�F�	���4x;[���?�o���V���lYV�RM'��R� Oŋhd��5�����`�q9�!f�{�D3X���Dj�۞�B�;��h��1�[	��_an�%����I;�$H	���@v�hd�u��1�n�� ���,�JιXx���q|��:d�=�c�4�k��E��xh{��Ii4��_'������c�V�4�k��y��1%x�R�r��-��<�X|��3�=�=nJsn�8�4�(�k��Z��@���:�� �/�A.����n�� sQ�� wī��@��
�6'Qˋ�f�q��Ͱt������=W�Ͱf,ы�����+ ��CN�Z���H�����]�@(��e�K8dd^�H�U�ա��8Q��\��ӐK�Qi�Ϊ�?T.�G��9��jόq����ZT�%k%�X��d�܀
\�-�<���=���x�BsEIo��TX��P����m;�F��G�(�JCξ��i��^!����us�O!+(Z���+���¤�"Z��d�dLÇּ���Z�/ߎɯN���d��!��=P={{����s�7���FK�h[M��d)I�ʋ���(�CˉMۋ���ov9S�n�"�-���1�䴱�x�D�'<P×�C�A~ �O��)M���wK�MR,�Op�AZD9�ޜ5�nK��h��0r�."��k��7ˍ����g2�x1e2U��NXa�<^�ǌ<����v��h��d#=@���bpu��0(ҥw�&'g�SZ��b8�Ma�)�7	~����*�L�s
�!�>ʂ�� �����}x�8����}7}���[$��5bD��R�%�}q|~����wMJ�NLn�x��}�K4�x��%T>t{���j^���g!
"[��v�����Q��2�뫆�!��� L�#�
�������Z�D�����C6�\:vxNE��o�4���=H9~��p�M[~�H\&qe�_d�I/�Nb_���l�)�*)5�P�,�W��M`?
�H<�bi[V<{`�	4�ʵS��f����n��PX�&η��͈�[�S�-�j�7Ec�s��B��=��P����������$"a��������hE�1u���o�/���������oo���&�do�Ji�D�7�i��Dt��
J9TJ��6F��}�캙�r.C˥�=rѴ�!���rX���-SFG�g���?��1*��D���f���0�݊@��1>���{�Τ�'���2�8�*ηy`l}�6�d(n�SpP&��W+M��S��tN*�� 9��a�;v]�7�)���*�/���~�;(���wގ��\̣I�2Ͽ�b��K+���y��HR?Q5O.�I�}���p�y}!�CH�H3����ԋ/8�D��+m�j3�tS�o�`گl������;��F����J������J��Ԁ�E����{,#'YD����