XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W]��J���
��+e�+��T0�gSEs�S�1l;� �B�����_Ͼ�\���i�Ѓ��dR_�h�Д9����Ⱦ�+��b��yUP�H�W�%��"�O����Z"@�!�k&�in$H�F�E�k-�R��<�%ޫw�ӏȹ���
��^�p;{ER	�by��,����I�8�D�h�k�66M��i>��k����7��rX%����}wE�b೚KF���Gu{/2t�`h�v2�Y�aEt4�"�9G�'��f���!�@�t}�y�e��k�C��2�xQ=��'�����q���Fg,z�t��v��J3Y�&�0�K}\s�x!GW�A���"<&�w��A�գ�����E�"�pڸt:b����bJ����5_C��*[�!R�&��DiT2��Э�8�;Ǌ��Ә����Ä�ڄ��8`X�,���6)U��YզkvB�1�п��qMi��O}��qO�+?S/Ƶcx��M��浫j�ftĴ<�a�T3Nr�1CF�٨,1�GS1`^`ۭ�l/-r�[�P�{�����8�Jx��y<��'@>��tyJ�8{����r�^�(qx^2�9��8onת� $������p<=�DV [F�����r�¥���`��ZZ���%�묳�`�Κ���
�=oQ�/�4t����'�:�������Q��-~D���O%LˇJn���ì��s��	+��j5q�U-3[��9�z�t�hy�D\��F�n�6������/���mᷬ~��XlxVHYEB    32c9     ea0�}�z�,k�&i�,��-[�\ͥs���L%�?�3�6�/��(C�b�{)�V-J�>�,rE�G+�m����7��=RF}�����ְ�%�����4������2Xڐ!b3��1#�fB�50r#�FW,;�5���%��E���WXe�}ڄ�>�(�/��^�<(�@�<D���j}l�Hk����8�f��zg�<'@͆]���m�&�~C#�S4�g~W;F�5?�T(�1�&������{��%�]o�B��{���>��M�XnVy�K�E���6�ƬD�7]P!�WJ�:|$����0�~R�A%k���^آ��$B�ͺ�YsAHS�SZwek�Z;�T�R�Jc����(����d��؍o^�
9�1L�G�Ƞ���+��8[]�)@K���W��7sɾwǢer�+�j��^_R��w�kVeM��`�~Q!��E'gmĴA�P'��U"n�L	ֵ���&��Te�d���*���]���cJAXBU�T���A)d���!9x�캹�Q@fP�+#��ujf�|���"Mh�EN,YCw�(�l#"c�Q�x��ՙ������#U�M��|޸v]O�����me��0���ީ��hR2��G��0�c�Nf>��q�eٙB(���tR�<��l�v�l\�H����"`Ђ%hq5JO�D��s��xZt-�d-'���a@:�E�q��`k<ؕ�\���Z��H�bb��$_k��z9G��3��O�*#X�J�.&�?�Pp"�{df ��9��<���_��K0w��ɤqed�됾��yц���j�~w�G�t�
�d�	~U����}�^���I��⧭�b �3Г�SO�˿L��i�B��)��]{���,mW�i? ��+.D��׹�!U;2�SF��9	̙���6�)��Pf�� UKz�@� �	f�5T����J�̀�#�I�}#��&�������HY�g! n]0�K�{֖�x;�B�o ��v�`{�J 	7�`i�X��u=-�@��l������(¤:�{g^ �@�"[�h��W=�Bۮ�1�^�I�*�L_>�`� &Zܒ�'��+ƶ<*U׃���g�������e�xx�G�Y�[�TY��ِT����@N9W�	,���)���>�l��Ƿ���B��M�� �V/j��(����0*�YŰ�n���51N�+\R_�F������%#���3�m3��� ��Ȉ��N�a��շ���QbÃ������F�w���ڱ�xqɦ��z����&���[�gͶ��6Q'eǺ`�L����Kv�a��,��	��ٶ���ː$ōy�  [�AFPCĮ]��Q�+��u����ap��@���o;Z���aq�����7��Q��b�U�dg�Dȕ�WQ�1`} 14ڱs���� K��K����w��P��D���ӹ��	%�n"]Qj[�WE//�pԸ�l��p��>��r��q��S�@���ǃ
�7�k~��i�	H�Q�nZ�B�;�M����2�N�'�4UK��P��'5�lP7���nH�5� ��ĭ쏝L��w� N����hU����歊�����܉����E���XRl�I�CV�'޹*�&����.�!����|3�����Qd,w�N�$�u��@�W��Z������p��r����!w'��7���<�9۶�X�b>x���U*.S��+�t��X�n��|�hXS�B�@;�t��Ph��e7�g��B\3�p�ʿ;�s�󅵳���.��a����#���U���$�f��4�]��vkJʭTP�	����nV�'8��-����&j�׮.J�~�t�ٷ�k���Ѫ��<ZkP����c���ᬩC�Zݼ��[�n�!?7��<x;@/�c��b��)����G����ɺ�H'����k�Et�a׉8 ��x)�\����1��Rh���3�`��O�5_n72�o)M?�S�wv\�{�#y%���t��HbJ���x�|TA���d1���z;�JD��1��作a�47�ZG3�O����lSm��	�����M�a�!�9��C.�*B��F�qc>w3^`Xp tC���J.S�,�Q�B/y5b���&�|�
��
)%��a �v�M=�&"XH�7 �����&�OV��d����2�~���^��y'�Q�x˟��|�}������5������*�U��4b�mn�����*��n�����Cx	�o8"�c�+�ۻv�J۰z��&�0�ƿ �9�LXc�S>���W�i�nM��4a�hU��z�y���ZBoL��18�k5�z�z�F���M���O3n
;}�`JJ	d��YǞ�E�	&5���
�S�L�������Ôo�}<^"��W]�"���5Rb �����S�����#Bsƻ~���I�*��^��sۛ�8H��>���(�s^���,��1��B?�T�M����Z{�����dE�2�ڨl�F���q?"f������ι��v�R����EhRNOA��@P��w���[1��qd~�K�ޒ��L{��m%J�
E.(��-Hl�<+�:?��,��Z�u]�O�-eP\Z��S�viQ�	1���Gy���##���v&x{���ni]���a�7��1��p��ɫ�x!_y��!�/wʥ���Hg� ��:F�?�i(��k=��}+R��sw�!&8Z�����k�y�予DfQp
k5�N�l��`���=o.�ȃ���aBQT	Ӌoɪ�-Tj�i{T �x�q��Ν�>�)���7�Od?�PwQ>Y�E���R�"�N��.:����Ս(q�]��Ǡ�ޏ��8�:��K�}�ѧ3��0��d����q��BFInb�c	qj�D��,�����#X��i@f�}�k��p�����x��+���%i:�А��&�в/
Q�%I�q�]�8�_/�|pTw$�\P,�S��37v7H�R�XIZ��Y)��[����ꀏ��_m��OV��6T�`�!��E'-��;;��˥拏Oվ��;�]`q��l��|	S����J�^���!x����-���?����;�"��Nsx�rgdvk+�k%m� 5�<@���oI��~���q��Y�Ol��Q�W���@f�J�g�t�r\�f�H@�A�n��1y�XwtH.$_��{xĨ�L�/�1B�c%�Wz]kav!��Nw�#9s< ���0s��<�и���#/$:�h�=�[���P�Ih��+�G����5x�k��q�nƫ9d-���B8�"񒪒[���+4�+�+5�IP�����1�M�:yp�Ji�W����̦*��^t��73�f�̣wu�.�B�;��T�bj�9�6Y"������>�������ԙ���C 6�5}�0�}Zf�e^��	1��5��%��pC�q��/?�!��/e�H����@�ʷ#�N��1�̊|�ק��|�
�>�m8�5#f�j�����;�OQ0�	�u�z�E����_���T^oO��g��+>~06]LͪV+VZx��t�Ƹ��i*��^����Ј����~Z��M�j� ���'���ϼ!_�����#���j*,��\l�^��;�N���S.��Ҋ<u!(�®��c�H�dL�4��E)]�x