XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r��I��h�$c7���j"�wz/�d UP�����pu���BEF��f��}	��u�?Z�U�Θ�?�1�*��M�Iu���	�0�s�!g4I��+an4rZ��&;��#��7u���᭶~l��]���7�U\����c4�`��� �a]
#�)=�������6l�cJb�XU]!�!튍KXeS���b]�[��l/ɱ�L�]��(H�ow9	׏]D\��)Q�}�E��eƣSԐţ7Uo�[(dP� ����F�:�=Y�{y���$XT/8)��"�z�1�zP+�6=��d��wv˥O�>9Vs���]�փ;!����O�#e�G�Čg�{���0�q�AxYomO���V�C}��'/�׻h����%��1F�Z<��oDri��J����K��1���X�F��~�B�.���'$��������+�$O|C�V�.��+�\x���.��y�$-���6��?
�X\�p�B�㋖�C8fȽ��:tLr��3#����E�Q6����)-��}ɠ����z��Lȿ��+L���#q���M�d����]��lZ��-'�8�f�p0`cD���gĮ,���ȋ�(��'��z~V�9���q�N��[�E͡�XӦyl�-���s�FMC�V��/�(�d�@��i��l��竦&��mQy��lt��{�N���T�"�<���#�^a��:ٛP��g�4�r0�>�� |.fĪ���7X�X�5�9���\`�V� ��ʘή�:Z�Y����(}�H�q=hXlxVHYEB    257f     bf0)�<.�dᲾ��aJv�K�Eqs4A�y��=�����$�5��&�T8:[@�.��³�S�V�'L�i# �w9p`�l�ց���8�#N8	dr�S�ߡ	6=g=����������0��kc7V7a����ʢ��!m�ye�(�6߻��>:��j�a;��*��}ؚ�	AZ^�c�Jgoo�F�{��z���tל�:�'�^���qgy���{�UN���J,�(Z�t�p9��X�Qq�uz^���+uQ��}���`�>Q�Aƶ�<�m� O��H����)@�'H���u͢8/�h;-ٔ\9؜��B����+ī��zQAz�x���hfs^�a���0�!Lo�,w��hƩ8ef�<^��O*M~g���1����N��I�OEel�;f���y:(k�&�\���5Y1ƫM�*�Vz�WƤͦ(��k8��� ��s��E.�>!�<@\�%�Ar�Kd)�n���fxm��Sf�1�-L<H1�$Z�'z.�{���U�~*�3������K0Z�P&�E��XQJ2���r\�O�����+�]<�vZe@�߹��,���-�Y|��{�n�?q�4}���� Z�^zm&R�=��!$��P�Uʬo���8>4	��8ϼ����v�lyj���h�'��7�}����FmsdsڅjYh뚡��3�6t��v�)T�⸖EAI���M9�"�-�`�{�W#
����{�	���ͭ��!�&og�V>���V�_+�N���p_�3h���G�G�������*�f���|a�h+>�v}|L��d��nte#Rx��� 
\��p�4
8{���cKf{h�/7z�2�i@��w��X�%�����mː�BS5=W�E�u���&�`�?=pۧ�ucM�W*�j5@O�Am�Gr�6t�8�F��r���ݚ�����y'�e��2V�5�=u �O�u�)�C�48(�M��@z��U�EC�W�����%�#HhGB`�T9݇�1 ����|��ީ��Sp!���\��KC��S�W>��z�� h��oc)���,oh0��R��A�rĵ�%�$o6o݇+j��M%e9v%�܇���l
�Nzc i�����^\�#YuQ�+�lm�|/	�y,����K>��M�vp�y:.�]D�7X0b����m�l��z炢k\���J;M�ל��P5���Ht�H��T�1W�ӊ�j���%"�����R�0����\��ٲe������Up���
8�F��ڵ��#���dYc��ۥDԗ��e�!-��>dQ�Q�=|=�s'�N~G�0�J�'�{���A����W3!/m|9���Ԃq���Em�w^�����t^�0��c�	�К����ǥpE�JɎދ���>� Οܐ��Hps;�g<z�<���<3υ��N	q��k^V]��̹�����9��^
]F��
��Գw�X��x\r[��L��:sf��ՉS�w�9�Hf-.���Kq�cu35��*���k2`��n��ϗI9�#DW.��o����g��} .XSg�C���)]#1�p�"� 4N�IC6sGy�]����C���±�xL�TLS�݁�؄�BV��B�a����!�e$��Ӭq�iS	�O�m�w&����{儐������{@<��������"�x*lO_�/,̆���i�K<�z=*�����ܐ+l�kvQ��D���H'��*F�#O���9%���{�W�J1�����n}a��2Hr�&��)��������`É�i8a4�}@t��J�yTP9���;���noH'
q�:��X��a ���V�-���c?����-�⛺��2�<�a��ʂ�6V�)���5c6������D	@��4S���f-����KN��4��Z0gC�8V�RGW���ɸ#eHf�,��/*?�e���îQ��o�����i՝��E�����5�
[q�j��ʉ�;�6�O3*>�ӭ�ʠ�m�=����2IuW��s��7�8�<V��.Mf2G�_�(�h�p��L���(E�������� ���?h`ﴯ���1"A~y�h�]��~%tQf�[z;���Ζ�ǁ��!3ȄP�q~�j�ih�"HBp��󕈁n�]����m�X�,�=������w(���S��E��ȒtD,��1z_ж }6U�w�G��C�-�+
�sv�lz�Ѽ����>���&Yis����v[/G��ze�B���7�"����<齎Li% �!��Ǟ�e�H�D�� L�d�A�h�Y��aJ���Z3�nI{�|��-�|eJᗣP̔V�B�Di��L|�(�����ڲ}�嘁$�:&}�#'�H�u�,!"��3}����گ=��zD�!)!q ���Ē��`]�T�Ӵ�- ���aW���ـ!ڄ,�zѼ�����qq�v�Ke�w���;W��M���J�B��׋��J��y��0'Ut��� �OR+З�km0��'�M˷�O�5��<2��ё����BeS��c��hQGtc�Ì@�wʤ����R�����M�m�:�v����3�j�H�	��ވ�3�'0J�/4��^�Gz3ͭ+"��V����H�M���C�����n9��A7��å�������g�6ڐORD�xOdl� �
���=�Hvn�%�<aq��嵏t��������^{ˣ%��e�2&�HC���`�9]24 [?��Ɣ����"��P#nу�<P���U�C���o�xc�Z�₯n�C*.��G�.�:^�#�=zXNWȤ�IP�@a�W����g7��k�\��gy*W��`��x+���1��ꍚ"I0��`�j����J)Nh��/&��f��"hS`����0Fk2îGz~f����՝ފ�c~_7zɼ�ᝣw]�6zIGP�.}���7!�!0Y{\ᷣ(*6��v��r����W�c>�R��+����w�lE ��7��k �}v��'tbl��+5u7�XV5f�� ��úe�*i�3��{̾��@���=)����9�x_�\�