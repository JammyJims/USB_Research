XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�z�L��/<<�2䂾�7,����dX�D
ٹt$����Y*l�M��=�a�Ϧ���|2~�����F[��p�N?=J#�8H%nk�O0�ᦆ��S�#g{p�6��>&���c𝹹` �X=d��#�����u�$5�T�z�m8��XCE�`�s|�IvL���NYvBβ{�(ٷ3��[���-�����nq�q�*�T�P0�Xuz�!��ǎ+�Qn�ȓ�	;�g���Tg���\M;*^u;΋X	.�д�>W"�:=ek���/v�+�&-$a]��m", P��/�v��L�Ao(�/&GTM<ߑ�oۇ �e��!'��U[ٙX��<��c�sn���?��D�ۙ�ö�]{���Ộ7�Y׀Zx��s��q��N�@}T�z���rl+���#�0��i�ޣ	��^e@�%�`̫�R�{ ��o+���^K�^���[�B����oq���;d5�:�}AW�%���Q�{7�
	��K���\�U�5���z%��SV5$�^[��eq��B���5��דUJ�\R�d/��j��k������G�$Q�7|]Y�pV���{P�Đ�r�ѣ��� �$v�ߎ5���ʅ*�'�1
;[G�[8_���}I���#A���+a�{<q��p�Z~�@PԷ���h�z����a��_�l�h��"���y���iy��p�;��w7u3�bԕ��w���>���^:��[��o%�ܛZ��ȕ)HW%W�?9�-�Mm��XlxVHYEB    11e8     770�.^q^��� &:e�h\�3�=�(����͔#�ȅ���2�W�d!v[���嚿�o��u�R}�:w"���pU�lR)�]_���F$���ʒiU�w���T�)��Ψ�!e�~7_H"Y0A�d��C4˴��(J�O�Zgؼ�o�>*}8��F(�H����v�R��+�S�R��T�@�GiT�L8���'͑{��� z�S(@Z�@�&DfS����ruG��#-�s�Ro|�w�"7p14��GV�� ݐ�����0KǇ�Ћ�D���"&��u��=��k�}Ѩd�;�?͍2l�s�9�C]��O:�7�ݑQ7ѐzy���hwr~R���X��v�_�'����ÚF+��'�W�_�}~j� �W�������Ყ���K�L�*'�KO�%�q�	]'��Q�,��"�M��U������kHʸ۟E�+1)�4up
{<%�*�`��p.$�Lu"\�V6��3;Or�M}�q�i~�<�͹�ð!�vKy�{2��܀�_W����/��}���޶����7w��r�|	C�S�'�C����SN�=R��#.%�#;�x5�%][(q��ۑ]#�h�)�e^�G����Z�%k�&gp���Q| q?U��]�G����N	��V:���'�kz�n��+�[���f�1e�@��M%���ի��K��n�
����x�`�g�9x�Lo�D�?�8�ս0�	c!~!LN�W�����a�1+�$z�nw�H�T�L� �/.@l	���U��7}���/�][j��ꆪV/���P/u�l�+����OQڞ��.Eԯ�(�{�U�ˣ,N�۷b�d�JAi�A�|xc�_��"��_z2WIĠ�3|
sS��O�
/�C�w��"��,˝���:�F6��o�&W&J�\4��^<�B4��&(}��<��2��N��E�����g�A��ƫo/���Qpǌ�ٟ��Q��b5A�[��~��KZ���'F(�)��i�.�����Xڋ�R����^��z��BV`�{]�/�	�tmx�Q�:�)�n)J���Q�,u/)��ḫ�=�6��uF3TQ�ls���4�NY}ɑ҆J���N;�Q$� !l���T�Og�&.���������a;v� b�[���l~KgB���ˎgc|aH���t;}Y�GJ�;��Puq�ǜ����}�K��}�6?�S=b��c85�nX�k�I�)�U���ij�*v�V�D'5�Fjr9dT�N��2�aC��}:F�����<9�s��sZ��ϝ~Y�<@߼�N�����ė2�Y��O��
p7'ɥ�<_��_r�:鍛L*Z���
��J��ؽ�S������v�-���c�Xl�t7�"-H������m�!��4r��bz���1� �!���^c�� $O�b$�9<����Mo��_���U�8M�S�F�XEG�����lSbd.AIL���q�o�ь�e�\���������f)�J�wf�Me��2�8�T�Qd-������������N�h�>�D�.coW^���m{'u�yl�h�OY�#��/�1�.c���7��o#�';5�-����;*uT��j�ź��̝"H>���tHln�-�b1�~B�ɼɡ����r���wk[���8���S^ׅ꤇�I���j����E�0�����<M�y��S�-�^Y�4��0E ����#ش��_S�-nw�Wh��F?Rq���5���faz@,�Rx��8ER��$�F�HS���]a�/q���P|�G1��IӲ�L����2���W�'*ݷp�%�`.�KX�L��4�I���u�"~ݖ�.�4�Y�o�0�X�6��H���͢t�X��x�ý�5]������֡����Y�x����'(��'S�