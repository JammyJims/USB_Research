XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o%�-}�ӭ9�3�	��ԁ�H*����<���u�:o�m_�:�őF���}��r�b+Nl�ݑ��i�><�'��ș��%�N�R17�m��[yb� D�N�H�o>�Ael0�Q� ���߉z���'v�[�5c��4��)
�*��8Z/��):����(�]8.�'��P���J�h��󉔒�'�׌|5��}bp4�J"���1�a۶��7`{���k��n���j!��'������17YR��V�-���4��P�]F�䇕�w���J���=k��L�����DW�W�#&(��5�o��DԵ �����ۄ%�r���ه^��p?C4m�Ǧa0i�Wu%�>3.!P$�2@<��9z�%�tGc|�X��x���*wצ��63��9!J=��H�\��>j0��U��;�)Ƭ�m�|C�ƃd����5���������I�7ϐ{]׹~n!�������`M����?���£-�7�=�G~���L�;[����� 8�4Uow`2�e��<	y�]�s%�v}���;�O	���.H��ⅈ�_K�0��W��+��,d{�\x	����K�f���{�?SV�)k"��X�O|���ry���Iॡ�3�O�6I�o���1X��=���wV��Ȼ!�2�U�@���˱�����s+�+�R�8�tџ1梍O�y���ЦI
�qe��m�nL�tq4v��XzO �3!�V�]o�ssu��V��$ϱն<�U�\dD̻�P�XlxVHYEB    507b    15f0}��4^-\_-��`�&�މ�q�&\���ģ�N���>�d���Kx�Y�0��'��|�;�oj5�7��O{㙏�`�(��1���I��q�T�,-$��R�L�S�V��. O<��36N��7����� Oa곯�J�*y���lò���]]�����a]�S�y�kFX �/AB��ó������4�Ƚd��������7��R����G²e8�K~@IY[��(r+�6V����D�8���_���<	�u��Ӹ�Lxq�:!U�b|F.6�w-Cs��V�9&X��Z� �3�����i��h諓���<5�Z�4�<U5��L�
JZ�N%����$o����Fwk��Fך<����N�g�Q,@?����F�8�o6��Iv�Pe�r�c�M���H���r�<�uyGɟ$ߺ��"����0�1�1�]�F�s)<☫2���=�&�J�b�$3*�vY��X�<�7X�j��"�d������()Xa�V��m�@M,�:?��"Jc�.n�x.��~�e���>�������|6M��jŉ�7�`ŧd.� |(e4��|�|��7p
ڸ����[@!뤼�c��R�UP[�w�pI`���nD��x16��,%���ee��㬃੔��������=nFeBj�G������Xw�¹�m��&s��;��tfa�j Ee��Q�,<P,ޥx�񪡱,~0Ǝ>vl\ϒ��]�*�E��Ӆ{�&J҇�cO�y�ǧ�:���`�h ϙ^y�>Xm�w�UXd⽓\�dUH����kh�,�v��j'A��Q�CY��'���|�X�_�~�F�u�XN��oDl"�g�,�Oa%��jb����h��s�ad��B�uk^.qH_���_ʺ�S�G�Ik
��m�'n��\�u2�p��D|�7�1$��h�a��R�]�7�(`��P��f�	�n5�r�Z��⍰s1����g��:L���"�	�B����,R:�qd��e���g���������(*�{D��`���G���x�Q���Ե���	z���Y��eڬ�� KX�����%Tfʙk���U��3�H�h�)j��4y�Ѯ^0E׃����%:j�1}�Xb��Q�n�>9S
�np�Q0��F�= s�E��'�6ŕU&{�@�:��aPFLU�h� n��sѕ��@�qK�]�L����h�$FuE_)\w��?4�5l�.��$i݌?"ᯉ�� N1�Cp��َ�rH�x.T|q~Z�b����o��} �,���JI}j|�3�*�hG4>7�T�L�~�?m��ٛ�X�#�O?��q��Ɏ3�E���"1�Qpe~�|���f��o�����G�
�M#<�)��O��T�RWBYr~Q�R�FBt�) �&7�`7�ʴ�%���83(6����h�4^�&�?ެ�*�%�	WS4�Me�Դ*O��R�����L�� ��U^���9'ҩϽ�w���,�H¯j��H���P�����e��5)U�a�r��Į��vm�iv�ڿ0#����4CS�����^�����O/k���NK�ôӗ��7>�g(J�*�^��z�X����\�I�1��>?UU��#�A��d���-�,�^�T��\�&�Vpj�@��V��%ĉ���|�#p;�?<�p3Q�Z����d��ܣu��1"=������B�� �_����ѥI���
t��q�W�Q�N'�mT��ay�PT�^5�*���o(́��r`��QkWЃv�㉛y� ��@H!�M���#�/
g?�^�irKq�e]o�5}�٢J�|a�x��R@B���L��3ܽ�8���{� �n)}՝�O�=;�ב�9/%�+�����X	�,V�,�oM(�v�PDHЖvu�^��ň���)����Mg���m�G������4�����m<����#��ˍ����N�n_$˥u�=,�#$\N���j��vD��(���k�so�[3
��k~��&瞛E]E2����%Ck���]�Lf�|T*�5�X@��z.����Wv9�ψ��S���{��V𧞓���0��D�V��zn�+�P��84=撚��7���ÜҾ|�P~F�a*�v�iL-̽��08y袎�C��W�mǻ��
�Ga�اk��u[�0��ȓ�>���E�qy&+QW˥�(&-�Ö�y���N�:��'�h%�<P����}`C��LS	���9Y�O�^uq�Jv���|�}[6���}Y}TIC6}��>��I��l=!��S�t�����-~�]��Av��S>Kw���^x�-۸a�� ƀT�ؙ2�棗ly����r*�����EҌyU�
��sq����O+I`J���A<���_��fU��9�y����9�,�dm/;��@��{%��[��l�^�QA9��.�~Y�QT2��z��!�T����d�0,)F#��)l��Ɩˇ�y��?��t��	��,�]ӏ/��,#���H���Ѿ�L�P�`
Ts���76�ކ=��̤\���(��:���^���<|A���RSK�����5X��<nX;�6L�����S~B�?��ҽ`:�Qq���{6;�	���n�m9�%շ�ⵘ��8���Ҿ�e�>Dl�,�L���ݐ�3)^{��)�a����u�����3FA�*�n�3��$j����t������Z��:��a;bIf��"w,��ddTZ�TiF����R�䝛	7e��%�q����͌ٚ�A^�K����/ymA&�y.۞�)�sɅ	A��0�<LI���B�� �\���5��Fw����<��ܞ��L�=��%����j��׍߲�&�TL�C�z���l�:0'/�	JD4������:#�HiQ�0��zXQ^C��Ҝ�u�m)1��L��G!J�W51��G"��)A����_��K�Kʖ�7�e��4Ѥ�l���}����BW �;��,�ұr�ĕ�B]K��:c��5|���y�B���~7�=t���^u��;x�vlA�y���ɡ�o,�&�hF��ƅ4f�O��i���~�+�-��7�vKq�Ap�K��T�v�W��P����O�&!���
~[�#U>`Ժu-e(vo8��L_���p������R�ZĥÆ)�bjzC���8�p�NE�}[<W��.<�J@�����{�=&�+��ge�B���UQ�*ߢ�W�3��h��Z��}^� 8ͥ�aӮ��[Eį�O�ר0S,�k�/2�8k���?�
$�G�-�J��Q�B��_g�aUE�����a���>z����)�����$�໡aJI�6�Z�SI�$�l�t)ت��u�1%�4���t�m�_�I<ǂ:'�T�-�GZEr�KЀ)���8��R,g"�	ĖZ*�Oߥb��kl��/"�� xx��oe�9ׂNС?&�o�=ӣҪϵ4n_��P���g��7��`c��w�.b�d�a��pH
����Ůa�D{R�3�T�k:���琗 �9/��e%W��Q� g�I7XUk2$*5�C�9�u�+�;^V�q?o���ϥ�Ђ���A|Xhf�������X7p��W���E�/%s��լ/N�0#��f��+"/Y��%����[w�Dl�/!N�y��aPS��,E�\����/��vGޔS݀��fN�̋k@֜;`>�*��}���LGCTP{z>�Z�Q9��N��x��6`n�
+�B��"���v+����7Hny�s��Eߛ��ZE`��Ro�S�٭��ZB�,����'0�n%r���`��jb�r���B%��I�Peg�@�U��|��3��i��)����8����i��󥂊��^Mu�j�'}%�R�	%�7MȤ쬺vJ��A�+�bӪѕ����x��1���mb� 
��%������q��9Fu)�T��9��9��!�����<I+8$�0��"� W���-��rn�;���&�o1����O䍁�7��eH���T�aͿ[ؤC^��[�E%��a���5�2���:%Uy�_n<E��U�����}?����B=FȈ��Ƚ;6�	����m�P%a��k�>�����,���w*��������;����p����:���@<9��#�-n�a��[[$�Qk�*8�%r����\ec��hO��Y���n��*e���ƕcn����B�n�6�D2�5�e��_u�j~J�O���Ÿ���}�y�i��Ś)D��\���my�CK�[ ���=�+�m@ů0�hd#s��S�yՀ�yE�M3��!ps�:Sy������&��@�X��.`��+(U����R����>��
՟��7O���NaOPN�^>�F�H1�F��8�
�k�������W���@\��a!��.��ΐ -��}����m�u�|��
`�_Mg��4_�W�B�DY���ɫp'jJ��E�f
�M���^����b9?�c�C�H�~an�Y�7�G""d�6��|F��{���ocw%X�ŋ��H�n��>$Q�ewS��7�G�����E-<��\����z���V���g#{��1zk�r@=]rPw�fR��d٧��Tֲ)���_���T_ޜ4yp6��"$XF�7H��c����
��n+��[ne�6��{,�87d-��BEu��'�� i�u���G�m��0�������L��S��r���0�dO��אM�_���"&�M�kg��޶i���2�{<Y�7�rU��>J����R����h����A�1�'�`sԧ��0 (��b����.�X¿�6,�� �;L����bl~�낸�"&����J;�m$g����"&�'֢}`�o?;�n��^��#����^�B�̹���P�	^��L	R�}�Ivpof��p:&��г���.��q�:"�����>mܺ�����0��%$�C�Xn��b^���H7E�k$7��x���=>��m^X�;���R��8�H%=�N{��O{�;�"~��.�b����>=���`�"øꑽ/6]�yle���l�p�-=�K���]� }.�<��m�}�Ib	T��7��.���6�����
	�w;�u����P%ͯ��Ѫ+Zң�� x�P�k� aΰ�o�TTر�^#˕\\y7�ǜ�Χ@*A�}48�G^��`��U�P[]�8*+|�񡴒-P�Ø5����z<�0�l!W�Qu�ף%��~��$=�.0wjˍ�Y��3�o�	I�p�B���7 ���0�a��YMeڟ�5Hs�d	zi��7P��M�/l���\�"��3F��=��cQL߄]X�Ӭ�K�JT�%��C������iɃ�\F��s:Ǔ���N�����!����D��v@��o��)'�����{�
�̏��q�D��	�i�p �������m��~�pė������cti܋�|���t�wʕ2���*r�6֫x�v�y,�z{P�n��ef��S����))�n��@6�X�*u#����YO��}K�Pq�5��a}�Ww��TY|.<��މz2�Q�譃��i���C��(��e~��.�<��