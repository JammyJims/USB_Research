XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M��C��輺�+N��1�6.qڥ�rV^�E����>[����M�CǚĀl���<^t�ڵӺ���\n��o[$4·f@Q�^�]��!��&,m����ic�<���z^��{��uHtۺ�𔒶n���#�޼M��Bn�4���z���u)īP.�Ж!*C`��t�u)�d%��P��:��gF�;[A�ϗҪ�VG��8I5�6@��٘}�!�o�fJ��u����K{�]�PgM��������&%զ��1�H���p�'"n�n�}�ԭ��ő�Evz#@׎�����t���$��ah�,y���'9R��"_$�V��B�.�=�ˮ0y�wa���Mg���9@�x�(�_]�{���*�<w�DB�r{�&j|��.o1O��v��+h��
��u�I&�y&�F����sI�=`:g�bq/aZ#��ޓ�����4��w���C�Z���<nAm���}.{�9Ny�=������.�������܅v59"K��My4M>�B:W����5|ձ�KfPu���AGR�� w��bc�ݎ�C/����`��ۓ��'.�"�����f�w��\O�me�>,p1��G�˴������y���?,�q���V���3��9R��q��b�}R<�K���0�5P���r2�-�m���2R����� :Ҵz�4'\�b�+N��Vjߒ�^��H3%��l�8���aiT��p^�R�Q�z'�ղSM�3��V;��-�*���ak���#&XlxVHYEB    1f0f     ae0���ۺ�]2�x�3��
Fo���i��r�}V�T���Jz|��"P�j2c�ඛ|��4g�^heK���î��V�ɧ�����KC1���:�^<
�m�*UZ�J2#Ѩ0j5����HD[0}&� \QI�pBU��[�j+�܅�;�>b�� "z�Q�a�v�S:]PP|�#�6��$��/�-`��q�QL�����̑D��S�ƒmcjd����� �8񲻈���������y�2?��{�ˀ�ͷ��mIp�k�/.�/��b­����/�ҷ�A�3<�H"��9�s���7b�K�dk��"�ħ?�yߣ�*ަ,:��Ro�x��Y��[�ӯj@��K����[�y�1�Po��3� �*��ٳi�t�V���u}.�5��
�W���JH/������S�E�oh١�t��|$"K0<�[³/�b�`��mUF��"B/�K2��a7��,�N#8H���m�|Ԟ"�����`R�L\�ܱ�!,߁�N1�f���u#�����>��&��^c�j����<V�~tn��F��V�����|�3
kOc���@ �(�f%o���/�D��(��*̾d�բ�:	��p�)�,��d�U>[�V�)�w�Q��FU��;
|\�O�>�Su��U�ޞz:/&�$�+���7���`4<�ɅJ	$�6|݊4�s�sC�/�2&����sxqN����q%m/f�V:�^d����ˮo��i��;>Q����^ 8^&����V�rZ�K���ɸ���X�A��2����";zm���2� F���_H��M5�ԓW�����r}7׻!�"�11�ݳt�7B;����}��2ׂD�ٕ�}%0 �oL��#pQ�~4�;?�*��v��.�]ݪu�G�Lk�>��+qq,��5���kKk� �ݻ��w�dCQ`˒)�VݨKּhJK!!u�]�}B��
^~xs��p���D7�FX{\x'&1�/�u��d	�c�\�xV�,�C�Bƙ5�$М8�ʄ.�$��Z߰��3��P�>��$K��g%�4��ᰔ�ޔm!�	���/d�~r�?�3v�{S�}��/OnJ���H���'�T\`��D���5�)�r˸K[Q�V�v0�����d�Q+a��M����r}���9l�:iV*��!�c�'��5얲y�8�e\ӣ�F'V���P�e|
�n�.OX���
0�ȸ����0Ov�Zd�0Gd�'����ڝ��P�n�Y��N�LR�(�P�%^���d�g�w��wݴ�S�w$g*���҆
ݰ3���p�e#�ò@�M��6ع���̇�O�������sP3nY5������;�L5�,uZ���g��W��JΘ�i�wa9}-��I��ܳ�9�P�/�F�x`P�x�&���01췤H��t3�:1�UW�¿gAI(Y�QN��+R�����)�g%^1�򌳰�(.������Tw��"E�����*>��昈G\mj*�����|�g��h	~V�pkU^�����i�t�3�a��v! �T9�g#�^�$�G׃m$����z
��[2�6)��Ȳ�4�k��帘SW4�U�U�[��?�y��^�0��EM����izZ��S_w��s��e�\��9=�Bb���ɇ��Ԉr ����F����ߦUzD"-��b��I\  �9�W���y���;��]���;Ɉ2;a"��0�"0l����5�����M_5�V�!!ed�YC�ʂ�N£33�!i��7�R����W���������oIȗ;��q��aT)��J�I�%>�I�F%�U��~#)B�h&���g��L��I2�`&�F�,�7�)׹9SP.��e�n�������)sS�IX̀��h��Y�̓To�o�f��_Yl����Yن�J�OEjʰ.�i��u�`��������i��	M��o����t��z�����;z9s(�P̆�W�Bx�
25�h���U��=[�l�(v�''Z�x ��m9�ׁ�Pv͛�m�E$90-��9��ݘc*&?�E��j�
�n]p��s���q�Y�����3];��1���}�
}�'=9��J�Y��1A���󳣏y'��@kAA��H�O&�*��p��䈨ԟ>8pj�7a�ޚm�~X�vm�+ʗL�:)6[��A� ����()wO���'��+����$��ACu\B����X���%�p��K
Y������S�3Z�ei�?�O�W���ZABȁ�T�@O��	��d/��L1��V�!�?�~��T�P�㾏��x9�䝂\��u��[���ό�hT�`����"�
���ļ�gq��.��4����pGvͼi�c=�2/����p ������ M(�!2��qKj�j�3��]�֯��͙��~V�k���8��눱�rtJ�#nl���ͽ��o���˧�!�/5a ã�B���Q{�c�^M(�Q���n�xة����g�->�D��]����� �{K�6S�8n)�Z���&��u9�}��ʆ������u2ԟ��L?2��{K?z�[� �f���k^6�-��,u���?��N�ƀ9�K�ʊ�S���(���,f�t�4d���������~���	�`1��Z����V�%䁱0y\� ��E|Q(ۤ��_�4�9ֻ�m�i��M��pN��3<v��81[���G�N�pW�N/��٭}x�����#% -`ub�j8a�=�&