XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z�t��3Z*��vW#JarI9��r���!�`e�U �܁$�w�p�����^�AM_w�a��1���	"=���*���q���L�w���ٟƈ��� KU}��BR�(��O��/�2��^��	퉅����T�1�fj޲��KMC��ʜ�RZM�-e_�g�}HE�+��
���R�g{��G�:�>�)K��S�S�7i�(�T�J�)L�����>�T}���#��<~n�
��.fS�i�V`a�B	��ܶ�R���B��`��,9��n���`����
���w��$>�5Ep��uθ�,@������S��hyY���3�@VoO�X�	�F�3֙K�Cf���S�6��2��nщ�
���
m݀����v<���p&*lt�:���2 c��i��g�+���(�>��ON����R�ڄ�l5��l�#���$�P
�V]�VZ�t>2�2��O�*�/�#�U�����'[���E1�N�nr����Z������������>z��e�(�A|ī��.]�,�}$��Iݯ�����,�G�:V�X����@��B�I]�U�:m���C��4.2������/��mTj�eS���޸r���@2��y��o�W·�zL����d�[����f��#�C���jf��;���\�q���֭��C'K��vYl�˨?%[Q�� �)%�m%f��F��k $Y��@�ֆ��'��"�����LU�I�e~Ϛ{>�BXlxVHYEB    fa00    2c30������^IQ6%��i*7�P76h�� �;�sK���x�]`�'h��Ԍ��m�X�,�x �"x��@�rUۯ�l
��)����e������������[�է�9���C���G��F�=9�&0'�[7��Fa�0�~�e��`�����:ٳ��`߭v ��îguJc��nY��wr�c|h
�Ofǹyڎ��Ӌ֛���Pƫ�r9�*�@����S�Ɗ�8�x�̫��C����3�6Y��gP�t9Q���Z,PNE��$�ޣN�^¥X&*����U�o�O1�߆o�PO��?��o�1@���r��r�p�,n��o'�����[��Eԅ��������'��ZԊ���%ۆ��:,TK��,� ���t ����P��
�'��T;w�o/�-߿C�_�⬶rH>�y\J�C	i��?�����O�X�y"��Ҏ5�$�c7�a_�h�(�I�  �?.�tM�Af�&���mق���Ǵ�j�����)j9�vvC�B�JȲ�r#;'M�![A=#>D�艧9��
�N�ɒb�!��+"g���*EuTRD"x�+5�T�}�2[��Cx�u��vT!�����VD'�%4W�ew��� 	b��UM���"tՅS��y	��r��G��1~d ��-��_�q��-� a.���2}�qE����u�o��d�����3�0ӊX�4]_�N��ׅ}���Ī5�Ǻ��7��A��4=�܆X�{��h}��p�W<:�EIs����h��ȴ?���O�[��^���`gy�;U 8�Biv�Ϣ����^Z����%�-a��Ӏ�I���&.��{��{��=ť�*/�|�R�+�:�ғ�, �(��5+@�U����$�T�-mLa��V������u�b ���6`w�!�� ���q��*c��c-PT�����Ǽ�CR�G;�b���' �\,�ʃ����A.��;�T'���2��� >����zF����KU��q�d��-��&�jUOg
P��7##��Y�ո�%�o���XDŎ�Vf�d6�Wߓ��7o��8&&����\Nlpas����@�!�j=J"�}��F��6X�2X�uJ�܅٤Yf��(䍁�
G��Y\��s	�)6G]C���+-��޴���5-,h�S�L3W��
��0\@�6� �萷l���n�����j���BS+F�"��q�7��0��&��O���O�#�P���s$R�E9�vD�N,H����3`0$8����F��!7�'�-M�	$�8CKڮ�Q�4"A��7������}��v\��b�p���୒y�'/�׺q�m$*d��e�����W�w�0J_�2vR��)2L��� H-8�9�	���t�~��0ħ��?�O��=r�}\��y�2�9j����[QY��*��ZcP�O�	0���"�|�%���X�K� ۧ�9m�?��	/up��*\��7��vl�YA���)ܧذ���qU�rN�)������vZ%��h����4ۀ���JN��Ǫ~�d�KNh�h.�d4�#�u V\w��L��������|���|T2Y1���:a,f��L���'��,4�ǫWv �'
3��s��]UE[�5����wf��-k�9:V(B,5h`Da�b�D�i��=�'
��� �r=��BʙhnN.Ȕ3R1T��'�l�"#c���5��֛�J�,H����b�&���|��#�}��>���,O"�	L�:b�W��m)�l:�����Nipu
%b����ʐ�bz�Is�7� o��,��}n5�!�h��|(@�%�B�/�<�{�	J���G���m��!�:�}&�s)+�E4ӅTQ="����
f�9�A��S�Ҷ[a���	sa��){>�b�,���Z���'4YO��J�ʟ0�s{2Or��o6����9�Z��]�,H!g+{��4qآ13z����lڋQ^���,�K�R�n5ɚ�U�!��4d�N�H,�WK3��v���?�ܳ��e��Or���Y��f�W���\4��wbWZ��}]��L\ģ���V����HF��'�r�4<��X-.�=,x�N>�&�嬯#/�V������P0*/����y�e㶆qW���{EՑ���l�a�&��e��>}�����%�V�s_��*RaF͊�f-���
E�ؔ�����g���hob��*6\y��,b�ȱ�tPأ��i=��uY��A�A�#��T��e���VmIE6��T_�{0&�[h�_P�J]�y�CM����EP#�sH?��=3����n �`�������ykf��ʎ��8di����9�� ��rF�����xh��ڢ~�Z�5�&]sP}��h��m	�GP�@O������P��O�Ǳ�R4E�п\7]�v��E�n|1ح�:��0 !���]_�m������>G=��P;�Nw�$wI�w��ɻ_bS�[C��� DW%��@�YZ6�i���BU���'ym��#W���Y�wS��.���A�U�����"�d��ZK��ت�th�K�N�[���h��!s�RT�yy����j��;���)�/��(��������q�1��V�T��x~]�(4~��o6o<F7�X �k�+\�˟9*B�����3�x_
ؒ�w���@��%Q!��-l>�2�#��^����h#ѩ����9�P�Vu���c�5Hn ?�����$����.}�6h�#Q$�OwC��*�����٭$�s,>������&6Jq̀�R)��(b�m�rrZ�z�#���	'����X����>��T��%7�;s��J��ғU�����Q�B�����"o@�^����iP���3;[��$�b"�͌}I���A��6�7��BE]e|M�h�$�-_cy���h��Cv?[����h���a����;�cz�_�E�	����*�R��$qa?���\�"R�PHh��
0B��M�3!�m��ZX�F5�9!Q w��V��p��,T\���O��5:_��%P�+�@�#�����Ԭ����yK�52�@f��'�d�2�� ,��h�S��_�ٵ�H�/��>��)�Ev �c*���U�u<��
�Ҭ�Tn�d�F��8^]�ͣ�n�<�B3]EN.�w-�����m�|�U�c�M�;������\rdn��V��!=�?�_o���K����M!��(�(KGp�vџh�u�S X�q`8O�zO����q�L�f��k�uRƼy��|�����b|"�{ XE��p���"՟vM���^fx�XI"�{p�@Tiԓq&r���]�8?��?����tO��ۮS��s�<]�.����mdK���z�s�G�+Q�Բ#>�e��)Pn6L�u�H���֖�s��Ɔ�d& "���	9���Z�b�m����R4ߞn�Q|(VN ��kgh��l�Sa6vo��rL]���������M�'liuTtܞ��sdS���=iP�`.�_@I�L�����K6���>�_� (/�=R�Ѥɣp�"�@��)����\��@utgI�b�ιO�U4!��J�m��Ɵ�S�W	��TO�\	��������2�&M͙�@��Nip��Ո�q��Ѣh7y�=�A��X����М��0u^.7��q48ǲ�W_��M�H�]<͞3�at�y ��"d�B���D�-���\Z�xK_k�l� YB��v⽊�+	��j�<k�
"���E�ff��9eQ��O�]hY��'��ӿ����еBS^��T�¦�����d��X�ǥX֢Sf���.xѹ.,#9Y��+�۲�8�D��>LY`yBse��IG��Z��0D+�!OD��Es�M�����t�#tjW����"d1|����y���R�5��N�x�Z�:���컆� li��f��=�l� �
�x&g�6o��h�&{��2q����O&�����K7���p�YOj�qa�@�����~$��sy$Y�~d�ԛ]ϲ�X�!�MN����墜0N�8�}���ay!\�HM�?b3��9������d{�<,��7i�!�]������JA��Y~���)�4V��y�*�y|�K��U�ͫ�R;�`��5~�/y�����,��#�!4�_$���Ko$p���r��r���[�w���n�G�jb��MQǻU�E%nݟ�#��s��Ԇ�%�x\2��	+�W�qw���4ؑ�)��V��aThAz��h�,u��v��M�����]�^��T��\�I63�^�\��Š����@��d���袱U�n̘�d��v���]�)�c�6O���³5�����v��
[��k1`���8�R�((Ss\��O"hw�smoV�1xF\A�Mn�Ei]f�9�^��*	�v$� )�'8nMB{-�m�P�Rp��yzS!�8M�8�_�jfF�p�R�/�[i�B�ߨ����4zvd�d��s��ȫ�h�'�6�l�Ih������th��A�������1�f?K�_���!M��4���?�exW�R��C�/"�>����N(p_�	���k,��qQ�g>:�7y U�SJ��#*t<9�eϏ�Ն<b���RE�n�Z)ͅ���$�\�����ѧ�|�h�h�FN��[9��d�y!�I�h[���Z����L�-�����6�k�|�<�����k�H��gL�ɷ�(go`Bx�0��W'��*|�s�w:�F �¤���"��@"V��iA�k:�`��������~t��X��p4�I��D�o��(�kGK���1������JZ��D.?|i�
@c����Sw�? ��D�h]��ҿ0F9I�$��UB�Q���t'c2�Ǔ7Syo���h�tL�͜�X�;���g��*+������.3��^�Ƃ�R���I�ғM�"�۪��z+]��O$��00�t�z��@g���PO���	�-濔_e���~�>>�̖���cw�<��n��<
�����t�{'^��3B;&�_��ׂ��e�Op�´���]rdGX4��L��b���c��4�٤ܿ�ob�h��#ɾ ������y���Pw���2����o��*�T�#���s6��m4���.Y֫$��y�L����֜f0u(2��ݽ
�u��,�����Ꙅ��F���"T��P3�Le�C�����:����,���w�ASS,��<�й�@F����Po����	+���t��Yua�W��>��
n���`�$����w
�U{�a�C�I	���h�����r���G	����|�Ez�W�
+���IM}�z��:��V:0zH�@��9+N:�]�T�E�����O���%tb�>h��9+��3����� ~��o�A.��`�	Q��E�2n�ى�!~D�s+�\r���⿓�?�0�V&tu�-<{��ە����H�7".^�O��@-�#�U�n�ט���'�%�+�0�������v�|�$�<Lڪ�ȳ����쌁��{E�ӌA�>;�&�L0�x*��cHױ���7T.����@ڮ�,we�I!`�%`҄!6����l�ͅ�O�^4��~����@<z_���ksȩ��g2�{����'�sj�m�և�-K;�R�_�fF��JͩCiD^���Ӑe�.YmI��z�CH��?,��+ͣ��?|x�begMХ�e�� =:��L�����ˎ��x���cR�bF-BHe����uy��h;T�y.`�+2@�F.�d4
�dȻY)|��� �Ϻ���6��߭��7b�Xصo��?�0&>f���~!ApdM_7A�lzjwT��
U��5�R���٩H���*����+�p�ܣ<n�����!�X���I��X�=�2��xnH���K���GJ�lSu�;��OsǅG�Bvk�U�s�4���jK�����qH��� F���)�8�9F��J�}�+\hi�E°�F:[�t/4Ė�GWJĵM�%�X���E�s�/e�ފ�q	M����J}��=�3��l�����Ԫ�W&�b��3puˬ	�0_��hі� 5�O�MI��ʥ�w�&1so0�J��cZ��(�2?���bX�0Ǧ��C*�N!/�h��^��k/���xh<�dR�Is	�`�{N=�Z��`xuV��>|6�U��x�
b��Vx���T�R��z[6DŢO�����-?�)�{��B'C(�,�ɃS<�c��J@P]�CW��.|HG'=�y�cE0p
yK;�7�K2��y]��$8cg���\�t���t�x"�2V��Q�KŊ�{���k��v��9����M�2�M�[[�:�c��v�Q�_���x.J�7j�J��	X!<#(�<)���"Ƿ��_9��zX��+���c�#�C�W���#�1�"J�����I��#�3x�h�_g�>�Ș���<�N�0{��!���Q�~;�{(b� �v�g7Y�~�ε�_@�@�и(�~����=8����E�д������s����/���M�67��8����n%�<0���4��U�7p�ˬ� �rW�iQ�YQ�P��W� ��^#�;�C����������^��ު4�n��);��bۓ#w/��FƦ�a\��U_.
;	l�:n��k�Z!Z�{��5��b�T��)��z�0_͙2z��z�3�룕��ܚ�vc�c8)ט�"+��r%~;!U�Q�|~#R�o�&���2��[{�"��`��W>�,oKU���R�n&a�<�0����|�le�.�w���4�~�w]d��J�y�ں_�?�ѥ�.��r�v	d)�⸾&��� ���a��ҵ�x�v�گ.�ǐ�`��N�)���KZ�����G��k�H��§J��*,����f���Q���El�^*��4����e�A���g���Ҥo0H����;����ey��w,Tx��k�����6�LO_��-��@�ɰ��+�$��[�տ�Mw�Q��
9�'��`�����!��։� xր�V���I��T=��C�k]�g�'��������O����#~������L#�*�ֱ4��S�Hl����V/؅��,�U ��3�3��G��_qM��f߹YΩ?��W�K�$�N-*$�<���F���@��N�tL�3(n�� �X`T|V������y�[#�l��A
�ǐ�u�z#bn(��vDG�I'grN����� }��Y2�ھE����#��3:z �{���tq�p��3�C&��{lj?��8��)!j�/lWq��t�����cwu<TV�2f����%Q�>g�u*�
s�C��|Ƣ=4��&�}�Kү��kzOOMt��1%��W��F!��YQ�暂~FthL9.d�	͑^d�� �;��w�-��[�7<����^ 5��xQ���a�w�X{��z7��#���}�<-���0CQ(�6(���yb�|󇐇����Ⱥju�%y�n��<v[X	������O��6�j�F�V�JC�vv���|��%��QD'Rw�$�qWq�}��ȏ���|jK U�qb��}���_��d�{f��n:���R��'�t+iX	H�2���φ[�D��ӻ�ݱ*/������9x�~���T[�3��E\h8_����r��@�3�) ���қ��AKbG7ہ!T`A�g|�*�ʷp���@s?}$k��c�PV�C�>B��"s k7�I~���z��oZ0HQ�P�)�aY-ڦ�P��G��o��#���j�˗V��hRjT�K�HRHT�W��Z�����:��P���8�H:F�[��m����kX�+JX�}��jb�|����Q�n��&R��p�s�3�]�Vn��y�ӗv�w�/.������sO��3 n���x�Ko�QVS� ��ߢC3^.��)3����T��P(�qщ�;=��9��g��¡��U4�b˵U`+w� ��4c<���5g��N��������..��&e�@h+@_P�����1�Q�s�I��I���"f=�;�� M�8��������}Kl]#�C��� ��%:����CeYl���(���.��$�4��[$����雃	��7m���AO���9�#h�	?􀗌�,�/g�� ��KF1��4�b,�D��k<�_k8w:�� 2�PoT�،��x�3�s�h�%)gIMX����l68�~�RCs��b|�1��7ȋfW�%aU�D��?�H�fκ,;���ukhɜ֜�ѡ��*����_N�k��b�m��b��)u�Q����>	�f���{#e�U"�6������=��u(ߵ�U;e�n';����+{�f���L�&��J;~Db洊\���~x^/�Hl��}��Ƞ"L5L#��^ly~���+aH��gd63����DX̃�ũ��^�]}�	�b�����;sK�4�hlJ���k_D�h�3vd#��B�x���g|֦�r�&M9y�\�௉vo����8��P(N�l����q;�����f�����0��yY���Cg�Gc�F_������f^}��ՒBD���ܝ��XS�#�$J��9�^�Ʉ��Z�&��~��ǫ��F��T�|�3��&�5����=�9/\T;�$�핖�3'���OI�!S��TW�?~#��Z��o�k�T�WT-��*�_�U�q����B������ab��b��k�,�wC�����ן6���*��[�J���;�~d��b�'�"���0<*����U�R��4���ʋ�S�W��\����\�̎���'CW���kAs���$.����_��W¦p�����lɖ���K~����jQ�;0D��)��������4��XY7�Y��b�qY�Ӑ&�8+&�������#&��?�}����y>�ͬt8R���|I�V:�S��� c�rr��{��� q�X�Χ��e���{��˚�t�.���7Z3�xl��F<Fl:�3L5� T������r��M��i���#�x͔x�)a�d�xr>G����v�l]%����;��SÛ�{�Il'�|�c|�;Ϋ_�����S�Au��R���N�s�zEfMjV�v�ۚ�óe�0�cʚjQܚ�Aʎ�)��?B���>�����@X��)?2�W)�q����(����G��R��A�Z�F�o����|�n��(��ìx������#�Zx����3b�T�f[���[�-��A#��
v
̈́"���d����P-����o&)��K�R���@��?*���ݢ�ɖ�AnG<�/\ԍ�1�x��mu�~��uo={r�.R�g��K!��']5Ϥk�-DW�WtSn�ƥ ky���XX�X��2����X<h�)5SM�F���9
��VXu��ja��M�����k}	���r~,��ĳĴ���ŋό	.��T(��L�E�M�ƝyC'Ģ��K��GP(���4񁖕D��o�ҵ"��Y�J
�cȗ�k��B
%"�
�M���{Hy���A8k���j�8��X~���68i�+��m��e�L�����N]/yRj ��x��%��U堘���;7qB�z��r�h����s����d���h�JQ�dm�FH�N��$��[�ǂT�� �;2��Ӝ,��3]�wc_�wN�Z�v_�Q�R@u�Y9C�{��@��N	m�z�Q�5T�� ��0��m.$�T��d̶A]�_��x��G�		�)�H�d9ă���5��U#�����
�iZ8<b��������|�I�����D
�9μ�o��'-�d�_��zrC�`��� l~����1
�b�MC\���&��Y$#áw.��5xTM�O �.��h�]S�
W��G1�H?�Y�AX��lI�}�>M��nL�4�7�̠�����\�/~`�}������8�!���m�+���5��B��鮺�<��c�\}��ڠ�9qb�{��ל��?Im�8��F�Wh&��Қǽ����2����n�ܠN���.L��ۑ���則�ɹ���ǦŃ&���^|��Lp����B��`,��@?�}��3M�ֲ�~��i�88�2	�l� �i��kN���NY�I�$�RvLp� D'И��2�*�g{��x;upy��(d�>v�L��m3U��Ӿ��iE_�'52]��/Є�1L5W��[��6����"ہ�� bo�_CïH��u�U����w#{ڀO�{���Ui�q٨���>��\>1��X����R�Ma[�R�]z�Ot6��� ��Z��=���1����A#D!2b4^ӸF�]���qjե�BkpeTt�7m8�Yz���а~׽�V�7��� ���׎wܫ��3:2c7��E��ycB<O�~kb�C��[�r,�sB�T �U�s� h�Dx���p�E���є3[��ϐ3����ҵ�y�Zj����E_3�PΥ&�1���$�7����Уp�RF�B�q�a�t����טԖ�fp�ʞ)�K������擄e��e|c�2������g�A6�Z�3u��4�L�ؕ}�evڛ�l�E�"�e��y"��Fȓ�����V`���B�_�e�4�Xc����ҬG��yY�_涋�I6�2��6tɐ5*{�m�}lW���G����|?�����`�4�A��Nq����K�w�_�S���é=a8�����G5���ʍ
rg����g|L���(�O!��]�׉�]0�5̩qRߵϯv�V�����c:�B�iA�861i?�}��X���p��y��G��$��b_I{u��Ieږ���A��t�bCT�j�zψ�Q�>�e��>� �4̺��tV����lnY#�=/ٲ�@�j5�B��&Y_6�s�0
�gP��.��g�8�"����cQo�Nˆbw:jd�����8���a(s��|�@y~ƕ���+�J9��-�Q��dP�1\�^S���_X� -lB?�:�tfUl�a���+u�ߍ@�8��:����-a(��I�b�9�7 �B��Ï�R�D�����/�:�qoq��H����ޗ�q�b�Kl!e��'	O�hoq���ʸ'��`H�t�s+��p>D��
���TO)���n����]O�3���H(�,Fz����7�)�)�TH���%(C^�0���H��XlxVHYEB    fa00    2f205�a�����u/Q���@i:1��ݰ�r�rrB*�Ԥ��m��'�vUd|nH ��`{����Ͼ�U�.�n�/fj�Q���D��#-��r_ޫ�Q8$E��(1��K����s[� 2�TXMp����h�]
J�f���ޗ_Z.+�� �����ÈC�N���(>���g�i}���c)�]��Zg�{cm:ydQ��Ƞ����K���������uNO�[�:X*�kHt$+�di��r!�L�!�4�k�2C/�
�M�~�iy�>rN Pf��?�tڕ$۷'�/!�O�;0_�Nz=��AN��Id8~`W!�� �u�S��{b���^��ư�Ƀ��-�!3;��9;/*��I�� �
۟�����uh��!;�3GK��2z�����n�6�j)��c��Aw�NʘM�ޝ���?��f��B����"���!���Lz��x�q��h���n���I�	tp���7��g��� ���1���^/
��jn��a$Fo�E���a�$oE�WN�JJL%dU�}<�5V��'͑F�M���!'E��ճ��z�̮~}���(EH��g;�$��O$��ϸ��Z\7e[�
ʹ�$��_X�ˬ�L(���ú	Ķ�t7?����*k��`"�N�1.�A�g�zݰ��n52�"�;��6C�q���>7^N��ϝ�������A��Q�>�4�,��l��椉fBzUl�� q`���3x��tjU�:��'��$�5�SP��i!#��K��iG����PQ�� �y{%T_Vy��h	D/�t��n�� m�H��q���R$S܊�]wT�.��3%�:�/������#��&�`�d[��{~]��,�L1@���ʒ�5���L?���k��x�{a02����҃�@?<u�Qa<c��cR�����/mf[J���!�`��T��e�~�?~����%~�XI�7�>��'��+�;�b�G�䜢����ܢ�����?u�n���\�u�a��{���v�B��{\��C5��}r�}����+����������c�%�6�Wf��o����}Q�'Սk�/���=��:Q��zA��ƚN-8w��y�a��u�-� �yy�tŬ��Y��_%��ت�J���C�t�ei�G�`ƚ�PѨ[b������Xjvz�Ȳ���t��p�����V.\S�lZBj�z�0q�jBKtoԪ��q 2�+)nT_��x�2@#�$�}�4h2��Ř��2�;p�V#Ɓ֨HZ�	���ڑY���{�����d��*�ꡆ
��/1��]F�c�iȩ��}B wv�M_��g�};��$U�!f�{`�	����7�A��Ұ���]O���S����O�l�)�4����z�t�[�ې�R+$�Sm�����ܣ�N���R�F"����&
���r�w����� ޞj��<�����!^}�Y�t�����J{�!.n	���'p�hP!�`�I���&1��=G9&pQi��=)����nM7�����@�R�5��p��ě!�|�����-TL?7hvVڈ6T{2�"\�>� �\�$X��V!���� ��u�;p�ܵ=#���Aw�u�cƇ�p�L|8k H2:���E�k�/�Um
�G)���P'���	�BN84\^b�w����o�KK��#�C!��`��Eq�JX��4�K1��Q�
xNo(ܻf�j�?��mJ$��uIh<�H7<g�ʨ\���{x�M�~�� "����7�e6
����mw�JC*	0n�S�q�xAC�o��� ��S<����ǲ��X����ģ����q��B�n1ꋻN_���X➹Z�~*�,M)�ԣWN �rdA�s��s�)B���;닩�l\�5���c.�Ħ���]`r��5eq�&	"�zܿXP>k�&߽���r�K�OsIz�^y�T->��t���q����&�#[W�9C���jO���-�4(���l�ڳF�/+�OP&Iߜ�vU!��FU%S#��6j�G�"���
�q����M�}qe܂�F���e�rT�	����N	B�#�xM��Z�LѶc�P�+g����K#*-�gכΰE�$��
�~�QK��
��C5t���(:��b�z�E��L�B�)3�$g�JY�S[|�EnڌZ���p��l�"�G������rx?�I&LX������CM_��]�Z�M�xLU��2�w�AY�����5�仾\��d4:�C ��S(=F"���B��S��_(���}al)�����	��8'eu�C�W�m:�/1�?�S���D�W�Z������~X���A�ɨ�4D�pd���É*����"	��d�<�d�N�Lr�S���&p�?��R�H����.�>K�ih��	����II���Eg��w�|\Q�*xq?�K�T;|�H�=���b*����k�ȶ���#v��|גM担Ht�	i�k���F\
/����+om<�ا�ᕧbh�`gl��2٪Qxp�E����&�T�H��K�[mt"��'����� |P#歌�����dn���,N�FT,�*Qc�sx���-�Fba�Q�.�����G��� ���s���6�?�Po�/��/��b��mj�h��M)-+:��9�7T��/	��(���q�E,4Ȩ�i�?D-6�K<�x��)�ti:U�-�k�3TG%���ܴ
�滚mi%����ʒq9�GmX����<!.���#X��E_C�	@뵍���d�,R�OI�%��ԩl�I�	q��b�4� ;��=��u�`�;�%��h�Bm�����]�3�37 ����}�,�,� {C����P��2 ��ک��B|<�FB��򢌇��7p��+��mV�H[GH]0Ơ&ւU��kwH�F�Q�@M�5NX�����l%�y9�>8"����w�DR��C�>Vbס�ڲy���sh������q�$�0��Y杢��{��@]ɪ���=�� ��q�0��ue+E����f��D���T�x[d�K���=���5�!��K���p�Țca#��Q(��z(7W�@��H�/��]~B�Xڇ�~���nƆ�ȸiM�~wZ���)y���?������	 �ѥ"m������J��ha��	T��),_�/ q*YL��s�~�:_?�4�ڨJ�M�j}D#��+�2�1��uD8��c(b\�Js������aEg�+���	�Y�*C���c�C��dJ�^����t`ԋ�L���|/h���Sv{3����x��a��+D	�)��TʛC+��5zF�.��������Դt�M�A����*|�/4�4&w�b�^�8V������}�zo���\��� ����_6���.����%��_�
���Η��#�k�)��(ҭ���c �85�a����lo޺�h �,�sΦ�r��W�� ��Yx�]��*�r��q�d���Qs(���!�����ݯ4�l$u�J�#���.r��
���k�˚�d�L\����;��~�oxj����W���-[����Gz)\�Q�C)�U�S+6)��%/>�WH{���I�+��<S:{4E��+� �$��
��:�oQ�e�?K���L<�|Lz��рG �����_G�sL�#k��vL��?�5����D�U���-��܁>q����2Dtf)1������n����*�ǀ���v9j��g�H�~�4����4;
��8_jJ�z�;�����#EL2�0_,���w��C�+�}�������7��M�4��cgXзQ�K~Ӽ���2f��D�H!-���*ߴt��x�����hb6SzT�z(a!o�bO��ز�U�9Q߰�a
����/�h[,M�!k���cn�k���Ev�j/8�掋�QY,]A�7׌�O��������Q���m{J-�A�ks�L�0�/��n�%+��n�eb���1o	�?�|�����B�k���K�$
�K'�y�J��Q�(  \A��_��`��j�Xo��7���z^#���?T�	A�"ɤ`C���g&��O���u"}n��m�0*߸���?%eF�s�L������ԓhWG����л��W?D'��b�תC�]�J�LT�W��.�*�_�����two=f�HO�L�V՞/ey�R�F�<�q7�(��E��k��{U}���n#^"!5;3��jI=�B�k�mY�1e�(h���Vk�
��Ȑ0Ox��/lg�d��<��Nm�kԸ��XC0���U�+�"�������E�
�Q1�)IV��"e��P��J��y6EM=��*|��m ���M� pTQ���t���G���a��),����Ă��>}gW *.P���{�_�=u�Qq���TW^�0�?�J��:I0�G׻i<�����|��&���ƞ��g� s@Gi�SC']���9�iX�=�"���F��i\2Z�-��Cn�h�K�Ne�3\�����~��j]���褱�	B�[�Uj<ь�αh���)�^�ƞ���n��sյ[I�_�No��a��!{@
�".Uy`����uPZuFd�2�߁���g�
��<��6B+�W����s���p䨘P���&��������H�K�e��B��L�A�Z/@}��01E:	t�u��f�������LRk;�a'�ty�o2Q�p��D�F4�x��5GZE��Ca�,.,�L��sM�oz�����ys��8s���sn\]�xD{T����/s����eP���"����ã%	�H&�tA�ك_�(�	�v5~���dy����ߏOj
�(x�=��$v�V-T����A�c��D1�>��Q�n3%`;:G��Z	��
@/�]#]�Om�Ä�B�}pr�5���)*\z. {�"(��rl�Pc�����D5�l����]�}ˈx��n>Ղ��9�J��*��
I�/���8x��5?��H�����ߣ84���Ve�}3��D@�}�ҥl;��  ���/6�B��!8�L,{�<��Ś�P7|�\R�>#�p���@�ÞW�E�u¶�:S �s{��rQ�7�-���2O���=5VR�>�-��>8�i�	�h���_��A;Q{b�̓g*)y�������v1,C*g��/�s��:��A)w�����V�3ԥ���0�f�R^�	��3�^���))�u�|�=�����v$H~�kF�Pz�h�L�:¤���$�CT�������L��e��W(ȥ��o���$��N�[t��ϞqsF���V�:EXP0�r١.qh:�en�d��XŤ�zfFc����O=.��ƮM�+-6�T=uyA�A�2 ѼK��S5�{q�r˛�jJ|�7E�{uKE�7��0��-�q!Ңo��@!�$��vI�o��/.����L���FhҒ�2ܭ}?��vwa�2� т��q�=Μ��Ը�b|.o�r_�����)#Oѡ�W����g����Ã��u~V6X�EK���J>�|��ub�U����u)Y���K��;-,�<bc�ZqK�̢xbQ�G4��'�`<��!/���~`#@�,8ė*���,Q��|l��4Ha~��g��}y�B�Ȣ	uI���*Z����t�p������Lf�k!���6߲4��t� �.�Z�<��\�^�
Th�%&%�Er�#D&;�)s+�$�Dl��!|�/�_�εy�&$���Թ�B�֪�nF+i�����Dz�'l��t��٤/!ب�:Fx�Ƙe}i��M�v��B�v)�0ķ;�����8=Bhd#sG)��R⤈��\�$0p�F#��$*��.R��؁����G@8�řPyb����E�ۛ�mN:E���Z�30(��V�@�5Z��'�؁;�c�޻�Y�dQZ�l�Q@�	C�
$���!����8��z����i~�7���*��C����}KXK��1�/�ێ���M\���$�ۦ�!�PDT���1诔]���y8<��M����Z`���O[IW&3��C��!�\��!��ϺH����E�5I*E3�ld�N<I��sΤ��+�Q�z��
_v��4�Fam	��&�� +��42���ݼS*�.Nwi�=��3���eY�V;�.Η�������K_ڬo>�u�Ǩ����n��h��#FF ~w�B`��j֫�M
�P����~'ݖ�V��J�����_�(w�h�
�I&ts��e#`/�񠬛F[�_5������Z�H��n�mvf�N6ӑn��m[��3Q�7'��N�V:o�o|u�� #}��y��$iN���|�	:����sN��u����'�h�&��wu��Ȕ�.��O�|�r��FI��)íd��{J�F��{�w1"�E'$u�ƭ�
���T���,O�9���ĵ������e�ty7�\�}��]��) R�|�j�4��i�hra,Z�-3E�e]��~���C�}��T�)n\�����!��������ѐŀ��x6jA*�a�$��b)� c>��E�p�kDF�@0�V�0�+Ղ�z)ʹJ,+-�N�������ȿ����s�9\�	.��{԰������.�)�C�rF6Hf^w�_���swgi�9$E\Yx;X������$��1y�e����i��ZNVZ��N�K�DU�;��g!9��M!V���e3>��<1�C�;�wA�9$�0���Lq��q�˿�jL�g��T ��	���e?�M�5�o��]	߂��pr%Ge���f��w$�`�\5�PRY8����8A�J�D��T1q�89n�U��v,.wu��>��ߝ� aoN��P� ׯVB����mz������p߸�l�	E��	k`��_�
�h
�Et�2du��Y��l~�O�m�����jv�2GJɮ8��\c����L�	4!Ӵ\�PKlաJ֡]�5.l���)k�0�u���(}�eϥ0�����m �so�U{��#Θ�������'I����;�{�C/��m��C�{.��&�,��	|��B��q}�f^���ʶ���5]���IJ
ɀ����J�2bޯMo������8̀����E�K��ۻwf�(mjbzg���^@qZc�g�����9]\��$�f[�`F�ki�S�9ZV�
��QU�v�%�K1j�Ba9Y�����.Y"ʩ��w�A���O����*]|�ۖ|��u5�cSW�Y�ǫ������۩���fa��j�����7mE{Ab����֮ۓH7�Z$�������� r%NP� 	fY�߱�$cI)4\�%@�꒯�΋�m��\w�R��0f�Ӊ��5O�C�!��|Э=��L*^u��5�x�̮�Ё��Q�h-����.I�xK�`��;�	-����3cg�_h�Rh"����lO�D4�HԐ�ۺF���[O���vtj}��e����z����*@���l9�]�l&�� �əN�5���	���>��{[v5�c��*^��YK��I3�^i|�:;V"�D�1�O���d����:�D�������|���1V�����472b� ��=0ݰ�F���νڵl'�.o��V��Z����|*t-:�'��Y�7o����N��q,���os���cI����Ԇ(]4ߞ ���F�i�}_��[���2�b�<�˛��	���{��E��j���a���l�*9���F�w$������l̑Y�o�Z՗���4Uiσ	N��
��>e��J��S��>�eՌ*�t(�a�a� i�{,�Iu�oC-�C�s��`�OF)��R o�B&��jǤM�L�b�<�KـS�A��Ħ�k?���r���USڶUN�X8��~�u�A��V>���T�l���q�c�x��|[{cZt�CU �ѷ�A�i�jG������X#];6}���8����7M�r�_�T�z�Xw�����,�˄�@�Ǫp��O�=�}J�B}4DNXrܸ<�y?~׉�2R)�yu4d��V�%�Dk>��v�?�wF�EYOҽ���#��Ug.�h?v/��P#&�]�F�}4Z x&KӦ�.i�c�}qKt2������CR�ܮ�j�2���6�X�G'�7�\�1�Ԝ؜�Ȍ��W�+�ۮE��n���rT���X�3'w?
4(��v���~�D�1��L�^q����������4��>7Ϋ>G)�)���c���q5s�z�xַ�EeUvŝ���J֯��ůi��*W�C[�����#�3�*�z�7��ː5�`�.��u�,�����$P�Ѹ�_
�լ�V�+\��ȕ&x�J�z�W�oK<���*�>u�Ks��wX�?��)������ª5_��%�\F��,�#`e�b��ڀ0��vy#�՛�]��;@JjUE��. �b�-�p�"�,A99���hk��ժ��zWh������/�L^#��mn���vY!����D!��]	���(|i�������l��1�xi&ɺք(�{�w:w��$1�oOَ
�t�Q�_�<�I�J���1Ie|ĉñ���������5!*_-�	�s�Ӫ����yλs��v��k�2P
~mO^i��H�Y���z ������F����<p�Eeҹb���u~tRxS��C�_�q
'!?c lt$0z�>K����p��U㗗�l����&��a8g��b�[H/������t��kQ	���Ϲ�w5����n>��^)C���G�h��EK@��4��	4|ep �z6�BJ0>m��li$A�\:)�����l}��WF���MtA�����%%W(��i��Y�����= ���	5�3��(����X�/��{>v������ػ5���(s��A}��TJw�@x1�D�r�Z�bH�c\m	�5���c�]�c��>�q����\��+ ��Į��hJo�Opy2=����^�pG{V����1�����JZ!w���t��+S��n�F?G�xO~���J�8:�"QQ�§��S��/"�1|�A�7#@�?q*�J2�3����N`$�۵� w.�U+��\l���͝� >п}���bV���W]6�^z!x��>���h(�����<�����j���؎Y6�2
�Y��\F��0��5$W&��E��U�k^@O$4���}Cf���O�6���,�LK?lܕ�z8���آ��i�(���L�f����̦�����ӓ�1�W�2�4������
~i�*�'c���! 虥�n=�Y����<T������)��	k��-�����*�Ģ�M��lf�F�_�r� j݈��tO9����0�(��b�%��u���DpW"Bm���u�b_�����l��W3���%f�|��p�e��fE��<��j�� ��Q�(���u�mj./�m���s��.i'�8��3�$�m��$��=L�`A���48�r%Y"إD��C�Պ�(������A��|V;t�h%�˨�\� l����k[M�Zb��^UL�_{/=��V�����.Ѽ�����*�&Z� ��~�_��O�޷��\58Q��`�"3V��-*�+�����)bɄ-�l�~$��j��@�Y� �,P�J������:�4�Q(��$/e�
�x�B�P� n�����KV�:��Y���2a3�"î���S��o�6/�����_�z6��ے`��怓QO����?��W�t��'���."�Ӎ����L�$&���a6ѱv���z�iD��U�̩���?Ǔ��d;D��b(���6���@��+�a�>H�	"Ɏ�],��S�|�ބD*N�a0��F��GI-�!��`;,�P�ΰ8sT�KU�
����e�7� ��nfU6W-!Tҽ���������
ɧ`����퐖�!)�7�ޠs�~ ���j�����|��^� �����"ݖ�U]Xu�����R���P-sU��`�=���z0�����#�\�7�샌��~����]?��I��B����0����u7pB��EC囚붺�By�PD�<�$�H�.��(� :�F�kNw��y\��!��F��J̅�m�-�o$Pt����[�~����X�]<ܸf��\�[��$O�TQ:t�}o�U{iT��֢ѼvJR
���Č����� ��~O�!t\�?H�[�q��u��J�f9��@�E��l2�?J'ML��ODꏋ�ח2�j<���$1(��ܚj�U�Q[t$�_��(cK&jj��
U�	����UEk[���{v"a�I�a����w�_f���CP�P ����f8[z۹UKm	\5|:���������y�.�`ī���7��Z\�A	��/&-���ʾ�M��.���S����@DX�����i�y��F}�3�ƿ��2�5�o�1�4�oS�)�[�l$�φ��4lU� �Mh�v�l��i�@K�jӘ��:Q	����2��VßI<@ ��碞��_�},�Ie�|M1���>�-���qkXj���L�Ҧ+s*�\�����݄��g�(�a-x�,:�g�W�af��Y1Ӝ��)�L�ٙ��H������6O��0�j�$�9Mz+��&��ӝ,A>�ˑQ�l|PKS�^ �\dr\ڭ�eٵl�BHZdaE��U'q������9��� d��t�[�	MVC��.9��"g��^�M����">D�R�yeu�i���5m���{C��"
/J������X`\[�F����[�&��j�#�k��*������C�l� �>d��M�:^�b/��"��(5b���u����Z��]>����(�m��7�E�H5@J]�,��,򄟍Gh���]{6�2F{�	�:Yb����X����lo���F_�S�A�?�HBp�]��Xw4��8`�E���<�ʭK;>C��j��a���x�T�FY6�Z+�� �����@s]g�
)�ͺ��<|4>l+�H���E�o�zoI�r:�Q��%��}�e�"cv$�)�b6��fD��
we#��2[�@���R�@���BBoa�Y�РIw�����f����n�V���~��˃Ew��p(��P�߻����k7W�oiN� 
 ����!x]/���Ӛ�D�Qs5��װ���D��sg9��dG�ȇ<�4gf��2�'a��xW�w��փ@��Q
�(Jj-�%ڀ��1�ep�M���r�T��}����U��Ϟ���Zd;6�ꖄS�/N��Ҿ�2f�7鬐\����-�ho;�f
ds��q>4O�^�M��}?S鰽_����^.0�Q	~�/g�?����Z+��s��ZJ������D�m�1X��X��+N����C)�\C�hK>�;��#�Z�<�1Q�r<��L ���J!�65x����D^�@��n���+=����K�c��<�P�Mü��y�|�e��O��$�6��������a6���˹�vΌd����m����;�6�����A[�ț| z�]&�R��\�~w�_m�ۺ Eyo�&�z�h��� k�Ĥ�崉xpJI.׾���y+�%C�7�;	��4�5�]?F$=��C֗Ux�%C��K�4ؤ���G#aw!f����,��й�5z���P��:j>A�x M�~��oͿݺ���h/��}㧎��k ����8�5���T�ح��������	0��4gST״�� ���RL~�`B�Q1ӽ�IsuyIQҽ�[�)]�F^+A[!;��/�Y���9��'v/��8eٚ��P������5���p��)Ki��8 �ꯀXlxVHYEB    7012    1530��$7[��j�˓ٝp-$O�	9�����P����#_
�����H9�X�D�2;��bje㢜U��~
��w���V( �E���?x�M:sx�/x X$�&m؁M�|�`�^���]2y�Ð�"ņ]K`�����v!fR�p)�Z�	dƬ�^H��O��������J�D!����m�;��2��le�� '��Cߐ��i�ڕn4S��{waàs��q�H^N�s�M�&�Nי�ZI�#}��@J՜�
�|�����g��+I��l�$EZ�"uk�0į�W�l�R��[HВX���˂��V�ش�] �cM6Y��Y��j���d�/A=�o����G����wOԧ�yN
E�K�ʠ')O����N����-�~TĹ��M��⠝�;�Os�՗�ϱ
z�g��q����
�r�9����KoKOCyrJ�J�/�e���8�Ov��Fd�/\eE����J�L���YfZ_��1=��v�U�IG(�68�x
V�?m��C\��q��2"�.V���5��B���c�O�bM�6��q����'��OI/�;_z0Wk̟�R#�	����f�U|v2n��r?�Er���Y�md��m��	�������Ψ7�\y�F��q�.]�9���fj9�<#@�}�*�K���R~ڪbY���0�5������d�X��r��tb��>k饊�����+��v���EU��p�:�����S<������=��
�wM��*T�b�5�����<�'�k>A�'L�/��:ջ `nN3��~��N$��xx'�ȵ-�m��׾�0���'� e�T��6Fy�� ,d��(��"�\����f��.vbV9����@�싛FƐ�q�+4R#�k�����C�DD�WG���8��1��x��jϔY�Dp8��_��[+��2��d��=	�gZ�,oE-d�v �D��&}���4�� Iv�T�ƚJ�o%<����M�U]����]oA򣠈����XH�ަ0�\yU���˰?�pI7΄�����H�f��XΈ�Ƨ���<���-�=�8*�GZ���Iq΅�k�{H��I�a���C�I�_TyZ�a؞i�c���+���6z���V���?P�O�+d���Sk�t��ѻ]:9��%b��5�չ�5��!Z���+HQ�����۲��**�5rI�5q�&�"a�pn�7G� �'^�T�nrb�D4D3G��#Y�=��pHe/�������@�a%v����ln��J�qǝ�҄�Ĭ\ 3���flA�wc���
Ѱ�wi�L�e�ֲ��t�B��c	��|>� Tŝ������'�����:+얥?;�8����s^��=_v��ծ�|, �y8���D7��΄�A?)�r����Z��(��*[o��uD�q���ߖ��p�8<�X��1L�`,�O�{��HBM�=��H?�Q���<����VZ�w����XP��ʄ�$O��M�j�#�~e��!G�p��3�+������ED���.g� �ա�
C�%��#���f�t^%{N
~��Xl!�nJ�� `���&�CV}���T�f贰��4/�_�����G�d���	�h����a�T�]2�5dĬNy������V��9�[��B�/���|� X��>�g���04H�1t>P�E��q����&֐��=�F��q���@i�)�U�b]X�+6n`WO޴t�'r����	;DzU�#���M���1�#Z�"�jݒ�p[S?즌��X9�E:xj'�ȗcc����~Қ���"9m�:�,���?/�BQ�ALH�Ƨ2ǯ+Z˥^�˒e��%��GP�0�e�~���9Һ�s6�y��݉+�1�e�� J�UiyD���SL�U��$��d@��*�:�|/CX[l�k���,��PQ|=A	���۪������}�Y�&̀�� ������m�!�r�t"4+xf�2A�Ȱ>+Q�:�u�S�����㧺��Ck7��Z�['�#n\C��xȧݒzQ�屆�k�!N�S���߆+��صP� "Q��r�!�{C��q��/tp��T�w=v��E���R)-d�.�ǫ��9���<!Zg)Q���4�K��l���.D�P<a���c��A�q���ڨ(e~�+ϩգ�N0h�3�s�z��;��2�tQ�V�ec�jt�2�h�����٫�]D���<���x�n����Yݬ���rG�*���%va@b���ik�P�<��������±�a�Gafj���B��fKPr�A}L>�+�7�(�O��	��~CЦvi��,��td����ݪ4^ȸ}��oY�*:�"E
-oAz�5�&k����
�p6R�=�T�	P�%�R��V=X�g`¥��夁��~S���X&��=��f�)&���/Z6�_�>��󵜩�����-ʥ��'�/8��hTi����)&��U!aU}�� ��o ,AO�H0$��F�:��f��o�n@���%,�%#i���l9b�E��ʹ����X�M@�N��qw�X�?���*�pt߼��Ӹ�o�}�7�_��&h�]ͻL��:���k5(ʵ8�Z٣4�ť	#9m{�������;˨�B�l�4z���/�Բ"A�N���G55�J�����.Ũn����7��]b��e��QߊT� �PE3���u�.���m�x_�.ǚj_��ۂ!��<`m�0p�<��\�3[�����p��?*|������p�n���pr[~�ɽ�no��'��|���0y �Y�rc���_���_�x*����4bM\m��I���q����K.Ho^�V�es��f��'p��ο��_ݤ(�kTjU� UP��.�^[{�
9�R2������A+`�M0�T��'I�+�/��*Tx:�)j��v7n3��(>u��Z��@2��(j%{+3�������4˪�jsQ�$��J�XP�X[S����=����X=qJ���yO��Th�a����F�x�B��4H���ڵ4U�
!�c���o^��x�Aɟ)+�?��o�\����)���OG�cgwh�b1Rw�/-j��`N̆�\aJ�CRޫ��Lo'� #���턗�D!�!�]�����rJ��A�E�/����s~��8��2�2���`��n$� jL��cOiQ$Lׄ:�ՅFuB�]��T���x�EЩ��T�3�Y�'������<���m�*coөn�´�v�/0X�^ ���t���Ʒ6�+�k��!�$�=�C%� ���d&H�D�X�h��'��K>Y�x?ժ�(-�#��;���:)�;V�5-�Y^�OJ����e������$#c#	!s�K���_�͉�3g��������X��/�eRq�
��`�4k�+��{�l�8u%��3^9�G0���	�,u\r��GN �Sg�d	��J��4y���Ke�LO��C��.��N��a/V乃�n��P�7�����C=�d��5wj��#<\���`(�mG���f����B�_�~��0@>�	�v����E]��o��%�e�T#z$cy-����iy�@n�}��o�E��Cq���{�fԍC��M:M��G+m4�`� \n�Vݙ�􊡖d��.�h(d�0f=�o���'��~�2xD��U�L�6vA��&k��8�e?�#HΥK��H=c�C���ׇ�QX���nm6��}I��M���{��U�NQ+!q�'�p�xa����o+O� �&��/�W��>�-�6���0��hS�)�hQ��t4��F�ص�KEus�SJ�9�x���~1|}|�(N��j&�%J)�7�hvMu�̇��x��m�j#��dy{�wTI�`��x�Y^d�`���S�g�Q����R��JC��eǙ
��Vɡ��#�ٰuװ���Y����p�u�py j�pq��r�1�I�<�BųZ��4��v��P�3f�L��B��lZ���L-����ؐͬP7ֽR�D4du�.��
�I6�̔�+��`^�V�����7��<�s��C��S�X2�O^�s�/����:��}�w�c����U\?*k�~�j�S^����v�lE��ɑ+��^T�Eg���'U�Ⱦ�P�+R�N��W`犹@G�1����#a�:K�Wx7Z�#���mR�u�]U_�-�m��9j5��래Qq�V����c s�Z����Y�����y���'r��Y�q|��<�nq�v���t�ƅ�߽'m�6���(F�+{/���3�k�(���_z�)��W
K����I5��������"�8,��8�kq|0F���a���H���/�g�4.��l�P��{
$j�������~���P��cqz��03:m1���h��
 tl"9��a��D�[�Z`�\q"آ[�uI�"�-��_�5��`يs�8�<Hd2���!._��Np�wUA:��̟@���"bԛMkD�R��CQ�Zm��pY��>��5��y��'\��o� �;�Z���K�Z�N�c�����ڣ���`�9����{���A��J���#2��3�=iλb����$MLX6Įl0N����n����떯>q��vUU?�����H	�� -���M�,w�Z��fâ37g+q{���h�b�+$����'C����M�߹#>�8��e/Ѽ��o*��0umPY-J'/>�^���sC��g���t����կS��c��v�{U�����������;�9���r<}�\���ud�|��q�P�1�|���{+u8Ŷ���}���\��:0�2�p`���u7�g(!�Ȅ��eE13?ʰ���O_�ؠP�]W���� 0�\�4\{�9.o���)؏���w�R�GvN�ʲ�0�W��w�"8���{�;�|%6�o/�vr^Kq�J E& �T�B�g0h�+��^�r�b
�&G��l�)��G��T��4ДfC5V:�׃����L���[%�;l���6z��F�[(�p�u[I��Ʋ��?��_�����i_r(��q[>St�-uQ�j,L�Z?���.=����G�O�^�n� �!x8�2�0tt���,��o>����.�w8�gjs@	^E_dC�����$b�X':[E�x��:�tx�T��e�]�.�a�S��}������e�5_��?Cc�b1�ԻT���9��"��e[b�5����Jb�h��x��:ǥm�6>�q����3R�&Ěǟ����'�AX�q���^��=%��N���B�s�m %�1O�l�[8z��J��5إ^��i�,���Is ~��;Q�v��&S�����df��zK����