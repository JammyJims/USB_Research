XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����9k~�J�~�^�<&V�]��wK��e����'��z$�Q�����f����^���M�(3=�0��(0Y!�C��q��d���w`g�_AZ9�M~�]/����R�����*��~�x���9V����K���k�ۍ�0��0;��{8u:9��
D�*�*-kN�]�D˭�X��Q+����֦h
fZ��F������f^&KUt��7B�^��t�9��J��@�C=5���bt�4� �\s�.���� }~�}���U#%��j��yT�0W.��}D�x2裑���ڞ�}�q�O��E[�EU^���"9Ú��ۋ(f	���)y~'�W�DY9B���V���Q\����z��$|�xtO���Q��\n���_��?O��9�@�cP�kƕ���У�X����y�yds꬧���_��P���Ԑ~��p��Z|��B*��@�AFp�%a��J�ve�Ns�4,��B� ��0������w���Q�H��ƞ-�	���_����-�*j�G�����y�Vu�ER�d�V����l\�����s�r�ъ_��J-��覶�I�R�z����-�2���dc�u�c��$�Y�?]?7�4yF6VIb*<4|�a�5���n�u>���f���ݻ�~l��d�2÷��]靨 ���MM$��&���x*L}�B�,�S�񩢃ix�#
�nؿ��T��2���1���d�r���m�+���M��u�k<}i+���Mb�XlxVHYEB    516c    1400��H���G�q��1�_.ٞ0]:N� �)�/�(��05'����؏� ����'�Q�L�3�C0�qZ�[{��̵��U#�{���b����B�Qg�$!m��[S4��LQu�OM���c;&�=�\�(iJ�a�g���ٳ�p�H�Ǐ��zϜ��#��ܥji�g�i|+�D��>�j)+���ON79��!��S�vX%:K�)DH~ F6��y�tW�.���� Ka��R�����o�yw�6B�y�?��n��9��e��:�K�b�������j���+s�	���^?g^�ǏZ:LU�|��qVG]�0M X�Ks��q���m������?�'+���Y`�&B��m�a��n��>�2G-B�I����.a<��k5��=��I[�����:/*��A�(���u �V~�n.���JtY�������v��;�'C�j��N�L��+���+R4j�!Z�f4�}��H�U�1�g%N�E��K����W��{p����l�=����b2-̋f��@������%�񱺜��D����|����j��x�" ���ܚ�����W���-X�0p��hvz����m�bw��p��M�kJ4������-�G�6�^�l�����w���ͭ�I~�72���\��|x'ѕ�q���=�*'�9^h�D���?+��K����O �4L�FsPً̘>@%��r���9�s�����dvB���Y#�u�c ���'1���Ԭ�"��+@ �s���K��z`���T����}�έ�]��}�ǲ�$��Kc��;	�/:��l>q�l�����׍��M�l��>�1�h�o`�-TT�Jp'"������Z{ ���rLXQ�T������=n�ށ\,r�˥!Ckv��]��;JN������\�"<:	�v�f��kmj�J���8��p�&yK��/�g&:̱d�N_E�R*���v���w��(����Vb���F���R0�շ��s�na�BO�����'AM᳭����k����]+�N:�H:��	`�xk���$y��fdjƱ��Y��ۑ��#�9'��o�^�[�3�i�Hv��� �F*�e4םQf`/`Ve�A�� l����c�K�m)I�8A����W8�C�8't��Wht`7�F��K��ݒQ�b��L��o � ������5���L�*�؏C��H^o�z,xB�ம���sE0���U�-�rD�\�����*�_��k��%���탻��>4�k�@L�S�S��p�<Ʈ�wr�ҕd�j|�fPvՇ��V2/(|�T��&'0y� Ӽ�4
��OV�Yta #z�QZ�(���w ��a'����>�5 �y�46L�9q�J�^5�4�|N�qǶ�Y�g��Ew����W�q���RC���F��Ĭ{���Kʔ٪�M��9c�V$k-��}��%��B�χ1u�/����j�σc)q�d�F�f��>���
��RWn��ݎ��I��J.>���Q9���.m���6��K~���c�}�u>���ߏ�ٛ�{�"��@1,)�]ׁ8�r�S��ݴ�����GSݍӏp���tf�(~U�0�#��q�V�y�c�d5˾d�_�(��n��)o�FAt�c^�~*�ѵk��7s,BO�������9��/# 9�Q�\=�,,���؏,K��Z}J��9>��bז.���u}�Hc�:R����CP��.d�{7���m�Ύ��`ڢ�h���q�j��̈́��1h�ո>zBZ�������ܤ���Ŀ+��q)n]��,,�R=|�g�e�_f��^J���Ae�f��!�h'��>�_��m�g˓����~R�n���H�7���9���c��i&!�::�u�%&�S'+�dd��H�R���a��>;�>���"���Fٕ��̡?%�+����Ǉ!
Ų�T%�{P�3%bh�aZ�,�斈E�����+�����s3�C���L��9��b�2�-������?X�d_x*\���=  �c2x��7���+�
���2# �k$���
���l\V��k��΋C+;�8�X����j���b�n`R�Sn�o�|��;\{x!`���u�)�2���Cq���k(�My����n�&�F⠋B
��_�R�ܲ�
5t�b�����:�u��S^�_1#h��Zq4� *j��:�4?hV����'�|��<}���1}��#7�n/�ݖp
i�$�"TciF��k6b�W�[?������]w܄`��0O�X�[.v�A�۾d�ϴ9U�e�.�fԯm�ʀ�1�4�u��Ǘ (����U��O�8\~���IFI�&C_]8k3	�-��ɀL���}�Y^�+����ͷ��7��^Cط��lʮs�l�c:Ӝ,��J�*��#���P؊4�iv�|�S>����Τ�<�P�F�(�=J����#��[n��(. �*�^��CU����z��q�h/mLr�"5�wo@,kE�vy��FS_f����ё'ͨG��W,`�����l2�����'��%�/�;Z�;��؅$ɢ�[�4��2.i��N4�dP�;�z�y4`�cM*�R��Q�ʓ�u�e��߹��iG�X��̘x�[$���J��L5�Ι��_!uy�f�G�|\\��y# ��2���b7���N���?��7�j�iF�x�j#��zS#���ȵ/#=�tj���u��+��}%�]�7�Δ�Q0�]��)��T�i�S�c��ڪ�Tt`|8Qm�+=�d���; ���*��%�Ӱ���M�H�6��n"��I���ᡥ�o*�ϟ?y.�,�󢶙|��[�AE�s��Fh�]J
As.�@@{��P���a�Q]چ��507Y�'t����I�%�@��w}������9f���?t`���<Kߣ��S�~���U�w�p��?�\ �.���:��<��0�$�ϖ}o� M������]?<��da��K&_=�PИ�H-�p Nkr�`�e��!�n��Y�k���@2�Z�)�B�}4�?$�E����U�XL�:���6F��?�_��pw\���֗���:|�iM{2�z�6h��?wWR����0�U�r������C˖Koo��*����enُ:m.%�U�qT��W4�����5��u�h�:ޙ5�5�>�$@92 ����{8�y=g����&8�f�;>p�h7�pv�҄�{0��������p��kXT��- >��I��FR�4۱��d$�ݙ�E!Us,��u��'OPy�n�[���CT��u�č
;_>����y�!�he%�<K�,es
������=��i��$�����,:#�§!�1��]��]��;��G�8"M`�
�EJ��55q��+�4�� �/�����O�!7`4�=̅�Ǯ5^�|��� ��|���gRK�U�9����Ai�d� ÓwH>c��c.Z���p�z��僢���m2N9�bjw�+�HM�V�55�w�Hl٥( 6��Qw�B:2݃9	e�	(:��:J�?I�����}.���6��~�9���\��b�Y�YQ�s:2vRJ`���kIXe�ff:Ec:�*�	b�h�D ~l����މ}_���&!��2�ap�5R�q$���D�z�T�D��U;��>1P�N��c�DV�ܙ�?p�z��W��y����X�-d(�6ov��|�����wRu6��$�����������d�ԣgrh�*��|��p/X�Ȳ	k(��R��4�,ұ^���*2�Lhg��8��>%��۽�ʐe.`�K���Z��i��,�;;*�+T�1[������n��
��͚Z[�F�R��t�y����ב��� ��S;<ˬv�����1���`�]�m�$�%��B���e� �,J����.�#��_����@FkP��<P������48�t�5i�o��{  ���j�7���lJ���aHP`;�rۨS2���P-�RR��j ���lH���h��Jk��\��������&�Rf`Z{�0��A�k_� ��-���ި���e����]r���)xZ��=xa�F7d�@ޘ�_� �4��J%_��j��3&�))9�/�Y�_��;�*�d��$6��i���!r�"��K���ӨD~��]�L��f�!�,^���و�b��K�����e�����&�/7PaI����SX=�#��n�h�2�@z�[�T\Bn���<�g�4���h���OA�7z|�>�+�;���D���E6��A�-�f�}�W,�qYҗ�^��`��ۭ�'�߽e�G���Ͼ��]�^P��(�Ƹ�|״1I+�}��9u�JT���1�y9��<�����$y�~���B��y�(%��� "e�|�\H<��<���^�b��� ��X��{����Y��S�(�<`'�)Cs�]a�B��q ������ޖ���8���,īlI��PX~�f�VC��D(�]�����z>���bɒ��-���%�;�ԉ2@��%�9|df���}M��f�@�XG��h�*͹�rAle~�t��t�J���r^�c�$��Pq��EF�]�kVoN���Xx7�wف�d��DX�>(��h�FX�J�����<����k�PƳ^�K��mƾ�jW=>ߚ��3�B��K!�Ϲ�t+�S�
<N�!_�z�-zW{�a�o�|���ܥzQ�C�`���Oy^�� �p�v�2Ny���'ٴ���,"�T̲�o%U�(�$&���)�2��c'8Z�!�!8���20��Ť��=[ۧU'l���	潌�%1շ��$�з���e�^����k#�O��B��2��	q���-�	t���P{���:�!
sB�~i�d�He���� _d�X�:=���.(_�4`���f�V�HW��џn�!ɁZ�6�~tOP���4��_���#�u�0�M��H��2�"�qe��~.��B�l�]�v�.���*Xi�t����<�<�X,��m�*�+��#+jA�[�q�r��P