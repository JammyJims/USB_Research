XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ZܺoKe�e������i2q�2Y��� @��Ŕ}���ڈ�,��-I��)b�s�A�["���X����K��p޶� ���7����Nz��ɴU���msJ��k� �Ύ�wt�g�)���J�ޯ��y�xxU�9�lmp<�M��}p�]���Ay	��R�[����j_��!!�0��݄_������.�ْ�g�6Uڡ:ҊIW[5��n	v!�?�D��l5[�,>bJ��y|X'�n�S�j���W��P�����W����ͷ�]��f���Egn���X���ԛU�1�,��H�dr��ټ�*ؓd@,&�+<�2��JF��`�8r�E��~/����*�#kj�ЇŞ�7���z*��p�{�h�G+�U���AIa����[D���x�������B���߹_�kcc�[�#˻��ep���Q�-D\S����)��v�7�5l I�={��>���	\�8
Gmu21.��E�Q����^����#���^IS34�r�=T$��kmW2���J�I��6�9.�yxb���H�K��z�.r��~b�=�pE{{̉���UyV���f�gG��OB^�OT����#�Ăį}��-S^|��$,`6��(�ݴ1�hV��0ˣ}{\ ���A1% #��U[P�_�no�lP@P�!��qˡ��	�-�V{u>2+��jhaR��0��~/E�}��yǓ��x�F5����Z����(x��r��k�nJ���یXlxVHYEB    57fd    1550�@��N��晹� #��q��N��1�%8������I���s�=@r��;��]�������>�ȁ�>�]ۃn�c�*���(��~�7�;�Mݲ{N��@����2�@�K���
��� �"M�ɐ���|��)qvv�wsR�s��&�@�=�T�i��r��o_��)�:Yb�Q�*,r$6ݓ�� ��(!�!�G	��m�l�gEi8M\
�|#��Κ�!�fr%1a���!��^��J��r|�r7A� D�P.�A�)F�ø�
��&X�l�`�aC�3���s�A��Bl����˪���\ ��dќ�!7K414ݾ7l��x	�ch�����;��pE���kKt �}&���^�e��=^�㠲�!,e��ާ�{#�w���^��KH�/��)�t��S$٣i|��%�-� �Q����3� �"�g�#Q^N�8��T�����W���US�jO�IrRv"�j<�Ҏ��h2���k�
ۥ^���t�B���B����!�{Z{�5,�Q�ɏ������8���S���{�^�[ �H����[��:�C����@�輽>�Y�LL��K�)���B�p����>�> D��hQݯb䤻�yy\	'9J��0;���_������ł�	��0+��]�7K�y�����]G��jV����\�:7w�h����8d�d�##c��
¯^},�w������ٻ�fG�_�,P�?��^��l�9��:��L}{��T����'�qzm�f39�*1�T��<H+Z��4��ޢIŌ�O.���G���o���H�U_7� ���Vcl��-:�ф�U_zm��<��tg�s�%����H{h���[�|M���>��\�����폔B��1��}��԰�w�Vj�E��;�������h��M��<r��0nDǐ�GIa�- ��u"�i&vH%8���&�({��ek����\���k�s�$2Cc9�Jg���9#�ɋp���}i��g��t9�i�,=:���3]е
��X�bg�z	�S�1%���{��ч����y��5g��٭��i�FU�*� �5�G��ߟ�9X���o(�;>�:���'���2���ؒ�۪�'3���2u��9q�/�8n���?������M�>��xg�3}Вc�&0�.K�\��4�>ᢥ�S�:=�+!<�����A#����\�{8�'DY��0vD�����)Ѯl>�{W�PH�Wע\��v%<�EI|�!6�Ϳ˪&hȮ�Gf��}0H��d5���ݕi�t9FU�)��l���5�'q<q��Nc)��ʝ��Wk?��z�F��mm�^��EԓZ���+Q�q�\2�Y��N��>�^���\w"����A^�v1�>F߃U�ԝ��TQN�St�N��Q�E�T�ڝ��;�5IߖvY��D��� �٫�P���]��?ѳ�.�^O2�N����:�٬�6��"��+�e�Q/K���1�n��])���0���V��Jhv���y;_DK��c����lpȭ�_c4X�o"V6���E��u+��'�Ks	f�ͥ}���Ĕ�O��\Q�X���3�l���OR����Mq �_ӹ�s��-��B�/�V7�t;�{�@�(�HH��+�Қ�2�DTx�
X'r9�&�f��ʖ#Zw��Ā��/u���gBM�1lؾ2�]x�IW������"P�Q՜�8�ES�����U^\��{W	x$!Ĕ߫v���8W�G��3u�8u�yE���T�?��������Ժ ��5Y��:7+�ؐ/*�t� �PDػ��{��TD0^�N�c�6`�z~����?l~��������x�8���q<[K�h��_�`)D�?�O1�Sr%<��>�p��$9� ��4�fU���1Oi�/ۆw����AXG=�J�Ϫ���AHNf�����/DdQw�E�I�/�6�<���m�"��a[��餪�5|�x&=ӹ
��d��UG��r�=�шoV����wR�2���1�䌱)���j��В��K�W[�����K�@�7��/[�!��dsa"�������R;�#�%`��GK���E�v=V���{@��aq%������7�-;��"���[��n��h&mZ�,;P]�1r޹M�;���S�^���x�:�
�S):w۳k,b8���g}�J3��CP�8�f�YbQ$V��I���{��^�6q)�i�q�g��h�vȣ�DHL8�Uo=P�C�5M(�C7�k-�]��k	{�\U�>��_K>�����ܮ��	G�q@�g3*�MN��B��m��65�ȉ%��ٙ:Z]�3@�g�e=T��iV�?G��[^��r50IC�M�%�syw���+��2>FhZ^`=^)x�M���D0�A��n� �������P�a?ǡ�j��O�X���)�
��8�i��EJ�n���c��Q��*��A��:���*&�:m�,���2?di�ĎR#H��,.�����I�5�F����4�]����=�B�EXA���[;�#JK���d��\�Tw�3'��,�M�!3��XDP3��l���t΍�����j���3�{NJ�"��V��@RP����֥,&���� %+�x�ƪ��E%8���n�o�1ףk��-���'���R���d�9�~�cǾ=�ȕ�:��S�T?�2i��~���n�sа�	.+ƪ^4g�:e�C�l�i֚�������7��4���x��c�k��&��d�͆G)�r�OI(D&��(K3�~=uJ�F_��]ڳ¿4�9?�����0�f4�K�]T"g0-�NS \d��ΐځ~�zY���̜��:�}7�l�U_�^���*G��xV��E���2��[���-{5�W�Q#n��_��H�<8.���pWqQ�[`drU/D�c�بY�<�I@���۩~�B��,6�v�m�/�G�>.���Q�N�����A�j/����/���l�V�P�Z��E'r���cQX���J$���8�'R�B"��!X0���g��D�n�킕4{���`�]�M��d���ͬ'y�є����px���7�=@>ɋ7N.K���������B��X��I�s ���,�XN���*L5^3�<M�|�!P!�W��c ����4�ָ!%Ip\J���ņ��b��&d|�a=1�~���q����҉��鴡2'Z��)��������SƘ?_�:���a���k��veh�\Tw$MA?s�פ	D��Byݗ����1�G:i���}�wa9=�
[��KH�~-.~�;��XՂиvk�9f�v�[�Қ#��K¶̠��N ��t���?0J�6��z�m3�"�8�t@:Z��/Y�����goR�
r]���6�{�TO��5o9z;Y�ehx�]�L�]�5³є��簸 }���]j	T���ۦO�q��o�@����Q�����0GB��X�h�O[C���o��u���)���X�7�"1��W�f4�&r��Q]r���{��XU 
Ď�D8�B�nxioJ~�'���Ǭ�xy��Qs�n��ęGޓ��qe��,P�h�������̺�<�ɣx�|Ylm���Y	��x����-�؞7� �O0�1��w��aQ�H���3��ގ��9�~�$'�I3��q�!�q�x� ;��BW";�Z�����uT4��2P�Z�{���dqmn�b'e5��N9�g�a��֡�\ʉ����6z+Q�5hQ�*bB~�.u����0�Q&@)L���;|2V�fQ�XD5��(�ŋ��I�&�h�Ńp���]�L-#sdL얃��t���;���tK�EYS'N�"��J��X���=���p䀬��.\˗	M:�=�����U �.K��O��W��o~:��#�:���(��?��h�q"� �|�'�B��g�u��v0;�ӿ�d���ɜ���Օ�0^~��WB;�ʗ���0�@����?�����/G������:R��g���r�=�+�p�h�uQcZqZ�-���+5�1��L�S�y���H?��W��ǥ,ۧ��#�`	=u�Ǔڙ^���*ܰ����
Ь�r�֮/s�o�zl�JI8\�6W��:�T��.��-���翕D���O���cxg /��]D�ĺ9fl��m0��?&�|]b�T���)��zTG"��6�8�,ѡ�by�M��
q��qJ����W�#����`��Ɂm��W�nG9~R�k7=�����d���=�Tly��B#��� ���`�*>�b�l������ڙ�}���.��f${)�| Wq��nk��mQ�C1��)����:7̸�O��z�;�n��`+?z�/p�6� ȧ��� |�ˋ��>��1՞ںQADy��GuoH�s������Bq�*��o�VRB-e����2�=*<�����u�=�a^�������\T��`�M�>)П�3Wˤ����i�DV7q��o�V�B����vz�|q�%c�lw����h���٘-�P���u#B�?�H�3@��FSŤ�����^�2<�����p��6�1#�;��KH�����Wk" Zp�\��yt4+��@ 9�g�}�����oC���-mmC{9�U'oR(��+�\|�h�}a��Z�� 3H�<�SB�9Y�-�bL���l��2������ R��հ���Æi�j1��k������X��/E�+@���	㉈�?P��J� �o����;|oQ��r���s��W�{�~��'��|�k��Ԋ��uF�Gl��k��
F�� X�5$�r�8��M^��wX��<����]�#鼙GVBAՃj.�t���1V��J�W��I$0��2@�%ez~f75ӟ7W��|���H
���b��i��y�ܭ����\����Z+}h׵��	��������ڸ��x�h���6r�k5<�vt� I�K�.��u���[}�;J�����^.~�Ɔ!�KzWA��R��*��9W�w+S�Ou��g��p���<Tu�w��v�!� � N�x(�P���'�	�qV!uE@y���N�O�{�wI{n.H%?�݋lÎ\S��"�I��L,Z;=����/�q;�O߃���}��h�=��%��D�`F#f<Ս�˷W��i�����^�ٙd�QF
X���������;����w�gF�:fT�2J��!�O���w���>|˿ť���.��6�Ϋ�''�\�'��{��7�LLh��V�.`�_�2�.�
���9'����a��{<�ׄ_��x��6��0d/�j}N�
��i�G1�B����&ί/����h��0a�nSRG)����^�*Ӊ��p���͙Ob�,'��Aj`