XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����"����	��.����-���d��L��f� ��]��C���p��&[�L�I��2v�O�W�r�9�S����1?��t�B��M|�΢5��At+���
���q�w�����?�ۋH�����+�����1{�%/�>��r���-7L��nCwJ�/���� ���Y�FcОn`	]�}IVk�y��:�O�<P��8Y֣鎿@�+���o+�O�Peq�1�jK-�C��W�Q�Df)BEr��"������؁��a�daW��1:�GUn�h��I��}�����������Q�cZ�H�Ә����=��� (�3*09o"�8����xov�(� �v-�|�����܏r@<�(�1�x2�7;1�T�������ހ&
l6aӧ�y��إNZ��19�7�J��(�ί:�H5��}��s����4R�<}��"D��!��Y�p�������+�V�^���>��@f��K?��@?U�H+��_��؊��ć���L�B�n�-\܎���{�c��HL�hGF��{���o��g ;U,���\,�%� ����ir�g��*w�@: ����z�rI�ըL��>-V,eæ�F�[�î���}6S�O�b���M�Q��=)>;����[��g�1)�+���7�Q��n��vXU��>ʲ�?�����W�J#��wh�r��=���drF!f��n�L�3ש�;�D ��jQ1܍(W�`�.4�W(�8� ������2I͓I�~�XlxVHYEB     8d9     2a0�p��Y��1h[,OB��#�y�h[����DnGW>�R/[�M5��r��8!��̲��F�.U佤X)�_��2rW_M�w�c||v��mq�`^�~k�Q����7�+�Y����W	<k�ؕ쯬n�9·>����	M6� h�3������{@��:�Y���]�c�a"9Ǝ��D�hR}_ܢ���ݡ�h��(e d �|Y���������>�#�<��j	l*{�|f�ϣ�4�ǌj�.��v�K$��e����U?�*��	Z�{�I���p�#��8,�i�����;�o,Q�_�Ob9g�z����x��Q���Vg;&gң?ĸH
��r%IX.��&3R�����w�O)�/7���9vʮ��12h�C8Y�/�߭�Z&���m��>��fE��X�52��l�<Nff�j���r`f����L�w�|F��6�PĲy����[��]Z%��5��l�Wx6H��:�l8
zNz���w���R^�����b��V<玿挳N��(㦋��)��U�l'_1���ds��ɕԿ-�����8����dj�Y�RE����"b83)�R3:���*<Z�CN�x�7F��l3�=�#����E��y���i�+_��\~
�t��l~���q�,~���i� ��p���s
 �N�