XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S�@Q�"����$�T���1�t�h���rx-�<� L�Z�S"C�K�_���f\�;�v�W4t�[�\����/�O�(�d~�e�91�6#����\)׺gcc�J��H9��V���]���5is��q��)	i`�j�d�3Z�G���e�`#��%(���j�v��qִ�]��H�0�wB�.��P�[p��i��v�|He��;�-Ԋ?����Rș5T6�'�Ǩ-�o�0�L��߶���C.q�`�J��dt��ۭ��'���裈��y�c ��~��C�o�ӭ�=dHy��1��ߪ��j��&q���P'0�q�6Q
�{��j�c����=M��7cq@��!9d�:hi�$��z�	Њ�yșƀ�_z���t��\�E�q��[ĉ��K�rN�ӊ~�0��F��{������_�@��Zc���7����`#�-�k�sЦ�> �,	,�]�\{Ѫ��ս�����z�8��z|�Ʀ�18ȝ|�O_/�5�b� M���}�㿟�/3��g"�ฤCm3�H��_�ذ�N�o�b��0Ie��S����mY*4e��\���y܊�X��XG/������3�o�:�_R"��R�+�n+��ʥ��I�R&�iX�q�R�Ck&��?������e3*��M�b��|54��.�
��:�u����Ԇ���2[a��XJ�L���ҥ�C@�f�\����4�cq&��Z��>4�����9�%�4 �@b(
6XlxVHYEB    39ca     db0G%cS෢e�	4�+�Q�A�&v��7��]�sU���1�B�GN~RyC�����i��T>%�%O�Q�����Ƶ҄��Ig��z�!lϓ\O_j۬Kָ�A�.H�>��H�=8^�@�*\E����hN�z��b��^8�ˤ��d��B ۜZk�����Y ��Č��m�6j �cj2k?۫��t���닖�~O	/!��~�4C[���R�qp��Bdh4�Y��A�?�<@'a��ct��V���{	b�O��8�b����/�NھbŤ�#���౤�[�}`�iTx5���lB{_LPaڲ�L�"�vC�:�k3��h�&v�U23���������Yl����lm�
�t͠��-���9��)T��|m�c{_����e�;�(F�X�#t8߀�;;袵��f���b�"�2�7~H�B}qv�H�����p�n	v˞s�5��;(����f&�y�э?�o&��n��H���6���e����'�`Yn�w�\J�M��`k�$%MƋi)B�̈́z�,��[�&A����"����P$�<�)��q�<�ӝpΊn>�r���ˑ����o6�S����=B��Ƽ}#�*��NE^.8 ;vTɖX�p�L~�y�J�4ԏ�N�Ln-���E����qx{;��s�Y�dU9�&�i\�np+UU:7�H��W����6/.چ�kg�E��G�B\;(7��{�v��(u�ђ�J�!h:H�!\��2�����+�ԣp�>�}`bc(�l����ec��܄����2��?�[@E�ٌ�֎���x�9ڕ�O`��p�z�����|�0�����Z�R5����t!^c�B4�hd�w���kR�0b>\��k[�S�������mK<�¬��^�üE���"O�j�di�1�P�/�_o�I����Bb�87��l#Ԅ�F�-�������������ǏXN���Y
������'M�.��{b�a��D�q2?�C2����t�z�'�g���ϥ�(�J�Ġ�r]��h3�y�J��v�����F���&qO���3U�=2���ɖ@q�j+�-l��3?oJ���҄4�����P�ՊI��R{����t���K{q�-C�}�z6;�~	-~X�B��[�쐟*L��V�i�v�Ԙ��K�%�� �Ym���~�/��xrc��v�) ��{D�os$C3�����F
�B���K��/�Rn_������ ��m�2���Be���YR��q���d g��ҝOӈ�E���� ֌K�^�I	^�]ݦ�x
�تy��q}��{u�\
���I^��k���.F�JJ�dG8��ӽ�$cQ��r�aׂ��N�����!GB�Y�톯����֔�幸��9F\�e�wT-�k�0/�P3��csS��d��y$og�Ղ~��@>k�$L�ybS�P��jR,����i��k�\�Y��.�7C]5n0SUoeҼW��"�x-��J~�+��Ȝ-XG��uyK&S���L�̶RU�)_���~�3��t��獉�nW��>�!�4�t�����H��쨊��8���X���M*<�Һ�*1i���y\�[�n�<(_�s��⫉3�/k��'ɺE��[�@�,��
�&��b�L	HiId��uS�}/-�i�m>bFH����3��[#����k�x/I5Be(�D�K�~�Z���i��S���W� ��|��(�o�zf���i[���d4(�8:Qz�l��@7=��Z�%_�|�XNa�2&���?�2�%��%!���{BӽT��\�4���d\	�P!>�,|_C�F��
���'�>�Q,�a47o���<Yjoq������vΫ�]��PC��,����ٱ��`�Դ�2)|���O�n��U��0?�����`�Q��JU�ܹ��rp%�?4��7z�e�n�"2��>C��y�bi��NE>c�-A���^�*�3��#�������ͯ)����_"����|��J��M�X�G�-L�_X�Y�؀̧}�۳���瘂.Xb�}�A�oA[e�-�_��dFXt��QB�i��`ҵ"`�P]ء�����?�m6�`i7���ge�T�x�"9��o{i����HN�ǃ�Ԧޣ}��M��q‚�C����1nᨈ�Y���S���MB� tk=;K���������0�}�ׁ�x�w�L�3>q�xC�k�Ѻ���@l� cx& 
H��{�R�Q�A�EW�����B�>�w-gE���+�E�ٹ�|<GLV�HJN]��e%��������{�;_hJ`��knC`4�ȵ��x0�ژ�/�M~��2�� JF�`V�<e��l�r�=��2P�'��SJ�"��ޒҁ&򗹪{ߤ����[X
��Yo�+��.B���X�6Ɓ�p�d%�����l	A����
������b��cK/܀v��+�����Q��u��Gp�L�������[�s���l�r1#ؘ�����i�=�qL�J(ۣZ�8]kx�2�s͵�Z׹���q�!F~�R�V�
<��k�^��ՀG���G��gB��Q���L�$#��pe	H��:B�@������.5��~1��@N)�f�����\dH4�(uۜ_�#�`��UD��\��!�����j�q����{ۑh�P�2�hs��W�]9�=��v��.�2E�6���J,鉰p�lsw܌rӝ�j9`�0@��4��'���g���G���O�t�]��'P�)N�KeXC���ڮEz%ޱ��A's��H���9K��O�sK�4�-yɡ�2�����E�iY�*���@�\�afx��m�A�,�]�l'���,�*��O�X�>ꖲ=l�>���C��4IDDZ����g�-�t�؎JҺ,�{��>uLșE�eVn���}�g	���н�x���j�^��-7���,~������.��^�-�N�r<ݡ�G����4(T
@�ty�B/�8�N�n=O�`���؊D0@&ń؆�-=[m�ɬ�^��F���X��oѓ�{���|��`|�A�n�)��%�����fg���,������g)Ă�s�X;�&���X,I��T_"���y!����~$�Aݶ'��o��iq��uE��rL��h;�_X�$�0q�,����I<}�p�xJkҩ���
���%�?U����ASj0=:�p��Sl�������w����fDn�{6i�U�:	Y=i�P�׷ Х�$iz,J(]'�e�B���xJ.����js~�k�%����H���kyx.N�����l����qS#�����%�U��6[�:���9�L�O���6}x��/3�GN��5_���P�d�!j¥|~�,k���.���z���p��F�r�Ih� �l�ǌc$�nLR�}����7�=��s�eMJ��P1Ky��Ƨ������xi����g���ҩ89��u7�]�ĭf��Z$"�