XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ܫ��?n~��e������3�`�I�x�x}p�UJ���rr���Vh^���2ᦅ��VI쾓|Ait{b�^��K�>`(�^ *�ǯf�k�����3aw V��"�x������ߔ`�Ǻ���+��o��uq#c��N���\#:��9���I7�iչ���*_%�/�����fH����R9����+ז9n^q��0��5�I1/��4~������bizv�H)�r�~P���cmEN[<�q�z�

�з������\����t<��� �=�6��x�9܍}=$n�|sg>�V9S�W���8_  `����W^h�i���8�%M�6���Ҳ:e���6�<�Y&���}�pDf�]q�:�7Th=��T���N��v�Q8��/�vT�m�-��& {"��üH�ѻ$
�Vf0��g
_;)dȲQK��.�^�����51�&d5������U�p�n�J��鴅�-�~�g6u����������a��͝���N�۲���|�-���eVt}���>r�*ioʂW��P�������,����G}����_o�������.U����x	�b��,�rg�l�u6����N��t���5�W�V�+�PO�
U�b&��WYl��d���+W����l�u<[ʊP�aʹ��반��a�<����l[�\s"���Q�؎d���3��<R2h5E��jR���n,2����E�mzf>C�B����}��As��G�7Xl��$��	XlxVHYEB    5128    14a0s�>.�'V�܅@emox��M�|AE��~MyD"H��g�Bњs �N1�B��
�;q;}�wS^�TJ��nwed�����������@�)�l�5>����WtW�C�a!��Ԝhhr��T�y�����_���|�x�ª�p����'<ds�l���;�%�u����/�f�j��RP��F��I�0�'�l��9�5	<��J�p��2Ui_KuA»��f�Q*�O��������@6?��z48A��G�K�8v������5����Y:���X��M��>��1ww��j-�a��}���C�uFi�a�+��.�����)���9P���QC	�ΔǴ�^��Kl�'�)}��/@H�|�(��Y�K��s.8sX+ZF�(��S@m0��� A���ݼ\t�g������K!(,W0�>z�"*l�����6g�Br�Yg�i	�w��`���-��""����e��#�u��0���Ի-_?gA��9�k��;�t� �@��xl*���e�wF��~��>2��_�LԿ�x�n<�vH��:�x&pۆ(2���˘��ǖ��޻_z�|��ۮ�����~&�;z�a��¨}������A�
�X�4"�Wx)7X�.��М��al��ǳ��!�*U3Ș;��v�B(�OJA��$���`�g�~�mt�&��!�����nYAVoW{H&��һ_cGވ�y�p�+�1%a�n�c��L�:n��K<�LGSyK�g��ϵ�f�wG6�ֈ�y2�RH���f�b���~�\�EL-�e�|�@�� N��t?P;G�;����� dj��C���q;�o��f��I��)=�,����%9���}��a�N��7�����R��r\��F@�����/�� �c���g�J��&x����L��W6e(�� ̒I���Ŷ*�pm�4h��>`*�q�U��Hz;\y$�,����Uщ�60qv�O~?A���Ԃ=Z,�C@�a�m��IT�2�0ݪ��=Ұ/N�/�l���u~�]��B Wʓ/[ZA6�R��Ǫ��I��<����^�(Ӆ�7�q~p��*>�����Ä|2��?F�57���`�9�Hq"LjF �8�G��v�=��FB��'@�O���ÐG��#eJ(�bݸ��?`�`tnL�p�d��yȃ�-�{:L��.��9��H� �f逴F'�Z�� W̫O{�<�b�Q]��Ke-m�l�(�����X��3:ږ<2�$Zjs}>��iw�f�Ǖ����y��&����6`����R�ެ<8���@�X�)��IR�Y]`lx}&U��2���#�X��1���J��*�']�Ѳ�}�W�c8kY��!�Z�z~	�Q�'�b��-���jV����i��TĨ9*����^9>�ˣ
Ҧ�D�3�[j�<6����7�k���.RN=^�-)��a�)֭w�q�Q�[�2��SH�52Y��x{�̳v,+1"e����^��ꧡ4'�i:2w*[|�<�d��!Ĵ��5��Ŵ>]�2	b�-@
j�>���*zj���e�:+���iS&�D�
�y���mJ�Fw����$r;�_��Bg�VLtM
�-:5^u�R��f&j�d�E�4c{�h^�^�?�5��c	0��S�Б��멣����?\�� 3�����R��Һi�g�Tp�%�
F�2���B�R!D�X�����]]v�[�t�N	
�>i���<��%����q�_�'���.n�l�	��f�01���2z����-]�:�ib�9��򋹉�ɜ_upT�E]#j����)K�ڨ>	��с9�^=��Sw^�(��71�.Y��<6u���	��|��K>0�Vw�i�q����%}I�	�o�Q}� (8�"ǢD��A�W��y����J)<a�D���'�zf��]b���7�(���@�dSq����r+���1�����J|Skc��>������˝�هc��ܕ� ���c]kO��c�:`H�!$�w>� to.���z�~'2���q���t6�`��2 蠟����
����.7��e��`�g����?���Q����?VH��C<�C�2D���T(��z�
�R�o?
!���G�8:^�]���y��������2t�|��=�Z�8�5bJ�Io8��*ʬ[q��rs1٩9�-Qe��y�uFD=e6�~�I_�J�<���,o�H@�~��,L��0])#r�� x�İ[�X3	��HRJb�%�� ���m�k���i�q��W-�5��x�!d�A�%�\��V�#_�sJ�˲D�r��蛔�n�qÝ�3nG�l@ϝ�3��O�Hδ)p�I��x��X�R���@�	��t��M'�A�`�YQK����G���'>�z -�]t���d�#w���x��.�.u`��&[<�V@�`J�̉lM�_��ʬ�g�r�}2�)c���ƾ��)ω����qY02v�;���Jv������[��6�͝�"�3nT���l�}ˢ���e]x�S&���&�@Q��.^	���a�:ڹ��~���I%�ژW���;э��\���IR�:=�8��-�,��,��F#������Xln/�}��  �R�e� Nc5?�J\)�v��Q�����L�^e�z`3��e@,T�e��S�:!��a�^ߏ����'?2Y�X��S�0 ���_B�z��+���h���a�l��gڜJ2T�� � 8-�/mEr�����4@Yp�$)V�$aF��cJS"�.��6�\��?��E�XG���K��.j�rd�q��)<�a��+�#��F���	�Ƅ��;�Ay~E�v�!)���]�pi[l{��`�}�dැO�{�9����3g6��e��dk4���&��-�q�F-�0�J˺rt�z�Ï"�nW���l2��Z�E෨�E��f���l���� N�>���&F|��GXyR�!��P�6uj\C��G�k�^IG;������U1F1���I�&M�wNS|$�j����ON��9J�+C�����
�Wځ�}#V:q/�ؽ�Y� ̋U�t��ĔF��:5�r+�J�V3�G�^��0��AM~|�ot!�T�)l�ӊm���0/:���D�1P�f|�1�u��Ԯ���0ldp�v�9v�� S�VPG�ET.��.y�����1�ܫ�<<��i-{�mk��E}o|3���q�g���������fNo����^ę)�,��>�i�[��w@G��X��$D��S�È�kT4�M���bHns��(�>�da���{2���!fr5 �,ǋ�;%�k2����'�GL�_~�.�yxx4�Y���xG��K�ܮ�D�k�z�{�cY�Ĝq�Qv4N�D>v%�P81�w�&�{�i����R�_�>�������0�:d�&�G{��ʄ�L�y��GC֊��0�^Qg����Q���{�!HmZ-�̛a���$����v:/Y��}��ȅ��ζ�&��{��<6YҎ}w�E޿J�o K���g�y�β�R҇L�����_'�n��S^���n���[��E�o;�^��Zځ-zq�hϙ%z0�jd�N�y�^e(	y����w���X����|C9-��:��������k+�b�H.v����H +VN<�6��d�qVF�=��Dӏ�:tk��R����#�pS��0@�+��,1 Kt�)	��W�A���9�`�Y��sێ@R ����8uo���0�����5��xs�wsj��c]�o�c���x�x�a���Q
o�u���)��o,覠�I��f@Rl���ټ�@�W|��OT	��V�<ثm5��e��������Y>j��u\�����>�B��^��>M��X�u')=���Ns�,��~L�gI0S���P=^�,#ٷ���%L �����/���np0I������6��t��$w:�Q#9��+I�ϴ��	�2_hVD�� �+V��[>/���卸�Q�A�c�؍�[�Cޭ/����SQ����t:z��� `�p�Ab� ����%� �3��j��K?���"�P���z�z�~'����%�6���궴σ�F��W��y	��?^�T�z��0I"615���.;�>��)m_7e���ɹ���܏��D�Fr��Q�����b��M�]O?����s ب�!�\�kD��g��;L��Xo��'��"焆���d87$K�1�������,�TdJ��|ZҪ�<�Pլ-�N{i����Cz�<����q���t��ÕPH�U��.���B�k�:��ꐩ�����y}r!�1�AD�����*qsJ�.�j���^8�97D�H*'�q�9��|���A=�J���75���I=�e|���O棬g�̨��]&�f ��x;N��>���zuѵ�Hz^ov�W��
6�r��I�����&�^]bݽRu3\���0՗�Lh  �n4khx6�NpGp�t*`���$t���/P�U�uW������tf��XJ*�;��n�i�ew
�1�3�����<�p��fb$&"U(��7LZ��i��j8	�*:皃�K���=e8J��5Įqޑ�	��Z�L�g���NATXvi��?@���|��L����F8Hڵ�V��M�*-`�k9Ps�g6�8 T�+]����;Z��ؒ���#�e��x�/���F�Ȏ`N~�>�3�RM�Рz� �VƷڹ"{������^�?k�� ;o�5�|���jzF��EMPo�?�8BN�	F�����h��A�D@�v�2�<pےBeȬ8�a5��H��\��o�9��et,z�!�h��;��%&_"���O0�R(�>�fS�ЫyƮ~�˸�(�	���q�~'O�m��IrT�1K%y��v��`v5ˈ\�������>������4ܦ;��f)������E ��x?��F���im@ʤS��jy���a�^pL�N�mz�}�[ˎ �r�-�ìoo���A�2�P��/�#���kQ󵉽���yt�>���ئ12B�b>EZ7f�UHa懷�rBd��
c欠S�����:(  �����P��R�bO ���Z���'X��,�o`�
g�\'�|{���ۤ �@{@����_q�w�wGJ�Y1d$�B�������gZ��J�ok�Lpg2��B RSӶ)�-wCNs�g��m����RߡTX�<~u�c��ڵ�� �@��tP�b�kZU�A(�����#d/]ڣ����s�g