XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p|��\��*�#ggj߲�/��[�/?����4����f�wn,.7�c����$�Y��\��+�`V�ݱ���gr
��z�Ӎ���-Z�y�x4�b�Sh^>�\�囯}��V�@�4c<|��<\s"��.U2j����/�<C�T`�ΰ(��<��Wo���tM�kg�@%����sF��y�j]�X۲*���'����e�c�l��N�
`��)MD�&��������%�ߕ"��͝����Ұ��ϐ�\.��oSh0iS��lԡ�{ڢ��Q4�n:�����*��tW�٬n�K����+�;�����Ml;�]'K�^��3�Z��ؤ����)���$g���A�uA"���څ�{�U	5���^ǒ��+oÀlr�X?Z>������#���s�j��+��Z�K�^4��6q��j� ��:Po[�w:J˾z}5u�|]H������Ar�1y~�%I>7+���I'���$�`w0A�Y����Te��fkp�n�w�<�xe��(���/�
Z��Y��1�v��㵭L	L0��o$C�s�����'(^v�\�隴������_� d�~��k�:IQ�dv��cS3+|�~;V6������O1��߯u������eI8}ck_�~Fq��e���mx�:�~���'�G��\6	m��((r�sA_6�v�5\�2�����'�B�9�
����d���8����n�(O�e	�4_�|��D�+l���.�/���ȇ3��?0�)�iL`�tXlxVHYEB     644     200� ~N�X�)�nm���Q�E� �Qvo\�Μ��u�10:c-Q�/�y��{�DN%�673� b��)�©�fj�<K�.�}�AQ�HJcfPs�LVvF�L�A�V���!$�F���@�*��W�u���%':R�{��q��3D�y`?����!<'�9����0��d�'��R�#3�Q}�;�Q!���7�s���s�sއ�|Uk5���E����ɇ谿�@� f�I=����X�-����3�t�g^��,	�6J
�'��?g�G�;c.Jj���&B�i^�T����`��gP�������˷�%��������<��zݻodw|��k�\a^c�+��H�x���� |Ndl�4����i�<�X�t��y��gf�z��,�bH�vR�F�M�f�S �N����_��Yk6ϥ�-7}Ԭ���zC�X�����^�핗�k�v�\��C�"�����v��D�Md�mP��6N��I�����q(�S�n�'