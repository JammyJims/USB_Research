XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� ���,�����wj "jG�2Y40��o7��\�W*#r���3���*��:�{�ǁ�xw�F-�Ê��?�(��E�,v�f8��F�[��.-��L��Z~TS=���-1��S�^��K��8ՒԾ����O��*�;>{��hb�u���Y:n]��&x�!V�b�T(��ќg�"�����G;�A�L��8JŐo�dJ|�(�f�<�z#Mi,1v�Q+~0BBY�|���ͬs��]U�ރ��v��}{l���w���#CL�&�p��B1��0
;�;�ʢ��S�9�e�۵V��~���D1�A׾v���R���S�@N���$y���N�T���c�h���0:
Ij�����e�i�'G�1�L��F�]U0
"��~ٖ-��ӷY���B���Q�(E�,��e.üy���ʙ7�C�������9�85���EE�4�;�}��	�}�������gE;J����j6�X����diM���+\�i�A��ZF�s�LO���آ�U�UA$����W�����_�,!���A�,��JȰ���j�����F��B75��!�#��k�b�ý��D��lc08���.�����܌A)�����nf4��伬	�����A�D��U�Ri�'"�S�	��+�5�2I��Ĥ+���m�3�^lY<8k�(�J*T������{}Ԝ\�>�~�N(��x�O~F��d�ԍ�w����)uw@z�j"���H�C5�=��s/I�QDQȓ��N94z�XlxVHYEB    482e     f70�D\f�˻�����OfR<[JC���e7�]�5�>�,��n:G5=��+-�L�S��r�Ǘ�dҽ������� ۏ%���f�7���Ћ��L>X*���s�SJWY���^��.��K������"

��0ܫk���Y&�Q�I���8�?�ϊh����2S�iəq��45�R�s9FOO3$��Vs?T
gTB������C�K�͡�]����)�p�_f�/N���a��"��ب�x��
��K��1�&�)w���
����D�F?���"��`����F�ts��;�U,M����L�]�U`�S�H[���|k�&���Q*�~ՒKF�^�RPc~�k n�8��X�}�n�O��h;��������y��B��.S�+#����Tj�dr�&�'f.#+ܮ.���n^�������\�zT_2�h��A���}rPtsn`����֐�*"1AU��}�kId9�b�U��c�8a7l�36($�h��������l�&3β��m�X���������ջ^���@��]�<��D�q�Uy��e�J.��
A���/�]�#��`Ͳv^WE$�*p�{���.r�&�:3����P��|�kp�K�7F�>��A��뽋�X��5�j*7�_1��5,и1�G�����wf�ƒ� �B5���W�VM��x��c��l�9�l�W�z�VT�Ru��hp�;���c<��Fl��t.oz�B_��]f�W\��ƹ��,�)§�{0�W��(����br��/���6���6�=��ljra4�9������{�@��P�i�q�S�`��	��}R���$���� ��z�M#$�� �GD?m7�Z����"P�bs�Oeh���g����k�)^� ��8��X��K�9�{w�<�Z�&&���q�9���;9��ve��/�$���e�YC����!3���U��`c���),�^�~�k�lj���	���/�����C|]g�-:4i��]�2��Ч�0�"8a!�-��dvlV0rL Gͬ}�dJ�[�o�`M#�/FUq:����
l���0~a�Y���&�.�v�fl����nF���`!{��[N�����A`(��n�F=�2�Ff�i�C��zY��J �S��ZN��&�z`�m�c����C���p��#�H���:��;g���n�S������`{�WI�^�X*���|<���o��ti�~9}E�@m ��;�O�U�K޵l�s�����^������jxxbyʑ��(�����<f���:	�%�W+�|"l�4tɪ�~k�ӊgP3�awӬ�#!|Y�h)A���n6��ɆKXm-��-�꼇���F�� ��W��
~�Q��Tb�Y�jm�3�;%��%-@x/IA��ͩ�\�yL�5�C% }���|" ���g�����fO@*�}p�)w�^�>��mZ\{!�o*��X%M��=��u�+��u$��j��Kz����/����굽Lw2��/@0�X;��@�-"y�:$S�P�
8৊I���޶څ�E=�G�h��]�������~�#˛����p��a�#�5w���ʸ��E0���@4{� -�������I�-�������@���}	E6�݄�
��~�o��N�ۍ��JL�%�iU�o�lP����Σ�O����<M{���_P
���tX�j.C�'5��f�]���a,��	n,�'_�#�f}���;]��TM^8�
/��_�Z.�\���ԗ��Ѕ������5HX��� 	y��a:�9�}��xl�&d�A�<�V��Z�2�x¨q}?=���4oQ�GC�dX�f�����XK�ƭ�㇎S�$����\"����m$���(~tG�W�.�|�K��K���Ŋ?��[� ��l�/۶�����9^3���ʎ�:��Z��6�X��T�</�'��?`����ڧ�����8Qg%y&�X=���sV�1��!������R�;�'�O��<B�Z����~z����p��QH,LE�*J{�3��](��5C��ի�ȓ��s)?����������>���-]�\+"�>�N�c�9(�?]�����2�1{�}�R���_[	�d��seᡢ�>(�:�� �B�q+2�`-��tE���)e�(�����Q�J'���$�+ʔ3㨩l���Z�z�g�L�-2�P��z���ziqg͓nS�Sr(�9�	��%���[~�L�R�&qqI[@m�Yv�?t0�Տ��S���%��tl�g�����e��O�/�!O�juiy���L�g'�i&_�`c��y��kV5��4Jǯ>�#M����*[o�l���?OC=�`"���}M=�c��O�>C">eV�b:�N�ix���bz�~���'�KAI�z�/~�J�fP�Q�Ka���]T=�U���H�������U	�K:/��9���2]��%E�If�ҍ���o��P�8��z��p���1
H��b��ZQu�s��]�Lx�I�/�B��D��?�tł-~��@��u����5,���m��[oS��{D�e[�N��NHݞG$zt�U�\��?Ӱ�)òٶ��y�t㲏U=/27�6/���Fϣ%�ms���e��������Q�[`F�$TVW���VA��yl���]N��C[m�T�,b�Q��6R�+��@��F�z3p�\N=��\��0��mZ\� k�'-�{�a^��]_�P�+�gS�0V�7�5T������{�"�ۀ`���\G}��(@	����
�k{��hU�xuc��胟�����=5�׹$�݈�{�̵����,'X�Fm&U�d]\��ldP��܍E�z��b�@*�ݟf�{����a&bH 	��,B��S�Q�*Ko[O
E�?	�<j3�M����^T��R׮ ������.q�У����o�	ў���c������a��z�Q�e7���p��W�s�F6��.r�t��ֳ���,��T�3dq�u'���4����M~M�z�Z�r�2���[�~�B/� ��A�lVrL��iî\\I��K����N��땣#֢
�nԒ����B�i&�!{c���SѨ����"�N4�㳁�2��T<�YRk�;��Ա�=P�}#k�%�����5��I�I��D������]N�_jo�D�4�b�Vx{���6'�8�i�'�ѨaE^�m�+����I!�K�;��p�cGG��&WW��s��P�J�(R9RS٦EӼ�.~j���
�ς}�!!<^Rc�u� y��0>�rЙ��(�Ccd���\4�Ö\�m*ܐ������_�5�p]:��}�j{dQ?���3/�2}���#���v�:�U����ѧ����	�Ѥ��Џ����4�"�:'ŀY�<��K�`6�H ��:���#P�&<��b]PV�n��0X�U��!�!�/DP���CƜP�ɨ�>6d��	��p9��A/�|_��T����>�I�i� 2GD)�Z�O�%����q�^T����̼���ʙ+��v�F����#4@�ei�}�3Ȓ�����樴Ke/h�Xf�J���]�ш:�28Q�w֞(�S*#u²������n�{�b�!������]���4Ᵽ�\���RÕ���F���q�F�����o�LܰK(��u��t��m�֏��~M��!�v�ss�<�|��Kg��Z�*���>��K��ÛbSŝ]��9YG���8�I�����겝F���5"1���t�\�.f؊(��k�i��"��ۣr�Pk$�F���KT�ۛDqt�1�:�3�+��;.g_˄�&�peG	�q�Fn�IU�lcAC��\}j.����ZT�����P�Ǌ[4<�rvCXs�j�^� ���1�G!y��ݭ