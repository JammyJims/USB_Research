XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�#=�̜�5��9��Z��g�܃7Y��(t;��ʿ�8����{(�2#w;H�ʭ�O� f��	W�J�b�R����֍�`�:�'lۖ�3N
2MA�X��R������a�R�̂G�����s��y�	&��
H
͔D�r��eG��R(x9�E���>��r{4�0�,�4�O���9�]����Gڋ��O9O�ɸb�6�@.����c��6�>�Oa���	>:�,j���ԁ Љ�,�<����ߓ]сG����`n��������D����2����]gN��C��lU�'|f�Wk0U��ȸ��)����]�R�ت��#�q��.��F(�u���7(�UZ��`4�Ebi|X7,^\Ӯ�U�ɖ�����5��bL+���pO��b��zHeK��n�7��ơy	��ڃf<�ς�����h� $�����w_\ �̀���fv9y<��e��y�
L��*'����������u�d�a��b�<��*xK*���{V��q֍rDOE\^��ib���Rt'|�a��[��A�,}����:�@�k�]����O�]ѾlE0��SpS1��$�}OG��e�]P!r�e!^�p��)Y����`X
0J)�Q:������@���H�L��Oňc�7\錣Dx�aX>Cs�u��Gl]y�*>�X�결P"(��:�x��ω�������[I%�`��������с�I})��9����c*RyJ%��l�-Z�zv��}\�c��qXlxVHYEB    fa00    3de0�@E��l������ތj%����Z��N'[�H�˗�c��	���z��o��UO`��v�.'�p�5��r�}-����|�Vo�?����L^LX��Av"�s��\1�n<�W���<���|)*��6�7ǰ@�?�.��j��T[kR���d0����Я�o�����IAcǑ�d��T���Z�yt�B��h��~����߾>�W| w��p�G$�]���~�Y�"�O):t{a�N�+C� R��i)��t�N��ܭ� ���X�Tl�o
�J�ea[z���X���Ͼ�܈��:rU�Rt�k�d�~����d �shi2Z�R���]A�M��M�_��G����P����$4����H��dQ�g�i37� .����j��@D�ʠ�N����i��D\L�ȋh������8����Sl�!a"���ڼSo��oHu�Ƭ�}��o�GK����U�6�2*���왷k�� �<��>H��Ѭ*)��t����q8�Ş�P_þ�����l<�g��W�#�|��[f�_�m�D/�8-p����G�Ub؆ڮ �2hE���9��ш�2�|t/T���@�ioS6� �j��bbt�v{dn]��mB��H���*�h����;���p��	�M���Fx5/������M����\;��Ukٺ�;�k0��{�b&�;��up@�rwup:Z|1+d<�!�]#��Tй`�����խ�C��l��V�P��}Z��e��V���𿨺#%穸k���i�d0����o�~և��
��f�1��@aS���	�jyо�=ˤ���ur�*����%�����|⒯]�Cf�;C���ϝ�;c�F�>�DҪU���;�N���$0l_�JGB_� I��o+���d��wn�Q8>іO�R��c;9���FA�����~���,�[d)\��T����\#��(�v�u��* ߭b����O7r�[22���y5ߠ�4�A��y$��	'����<�A�$6��0��yoD���J,�������E�?B���k�[ib�qy�U�bߞ@ld�-/ɍp�)�#�N�)�$���OH룘���A�i�LC��
i�]�g2������� ��C���A�g�H��F�m��;57;N��l���+��.��Ϟ�gI��v�u<���5�E�9M\��7<�At ����C� �Ԭ�j&�m���.k��*��h��?	� Ck����{��
���qpS��Z
��6��B��1��l�h���L,p���7�<���FNe?<b ٹ�?_{��VZ��`�k0Bh�'O�Q	<�ݖ� ��<7e�Y�l+���4��b�[]��]�*bCX@����M^E�x#��_�9G���D>C�1\u�n���#�����b��9�8�C�j��K�?��Ϲ)�/u*$�R��3�s�	�3�u�a�у�r<���`��㦫����p���Zc�žL�P�����#Kusi��m/|���U�������ˤ�(�W}$��+1�YӬ��+��N+�kW�w�u���:�,��b�œ�}�	f�=A��.jR�uf�O��X��X����X�캟��n��~���c��z��!����@�~�K�]>뚽H������1ˍj�`������k�Ȗ%�F^��,`.�U�|�Sdn�����)���n�J�}f�{]����_tSFi'5��L��ږێ�C��2�T�@�k��o�N����C����F�cᔍ&�J�4�b�g��1%� sY֡�1��b/�����<"�����d@r����.��K��_!��J�z�{.�;��_������ڷ�&�O��p�&���8���a���B6B�9߆V�u+a�ȳ��,?1k��e�}�g.~]>����m&ݔ��ij�o��~��,�do/�Ӝ��Q�B ��&p�ex{O����qv3��P?�cɀ������B�{#�crl9���z"9�i,=22L�8�*d��HbT���L����?{M�;k��Ff��g���{Q��@����]9�J9�#��T!�ዣ{���D��I͵z�h=Ӈ;��Ȼ��7.���E�5�j��y�:����OA��`IHS���kl/J����)����DVU�ܫ���u�b=�T��{b�>����f��4LڗM����jD���n�^!�l�<{��nk����ƾ��@Be�][�
^G�`��"V߰�k�n
Y�aG6H��ȝ���,����w��̙�Xɢa�Ze��˭.��^B<'�AtC�dw$+��/k+0%�9��H���ϐ�%n���]7oæ@��;d�g��Ɇ�8Uú���m�v^1�s���de�_N�
�6�w5��|D��4w3	��l��Af1|SyYQ��5�m�4�!P�PA�G��1Mej?���V�&����q�摰���k�`'���(Ł`�]3�,8��r�����	'��:�9Id�g�����4PO���c�*�0)&V�c[�ªJp����4X-ri��0j�>:�������To+�@I⃉�k�����#P�ճf����t%��%�R:��e��s8s�'�wf 2
�FO���o��S$Y1$��N��,a*�Z
c!�N:�q@r�W�U��V�ד�X��ҹU^�ܖM��6�ǽ���XCC�e:g ;�3��g\�^��"�M�5,+��0��P߶!���GQ�}Xr�1�mX�J�3>A|�Аt&:B_g�1=JN'�ބ�p�!Ku���ٖH|b%K��Q����C�M��$;ڪ�:`�-%������i���S��>P�(�,A����ᥝ��+W(4]�]��HQ<�n6���˴=�Թsj݀@M�)`���B��fq�T�D������ՐR����Wr�c���qoV��8aL��p?G�T�o��_:��0�� ;�F"�?*�J�3�7H�N�3���(��Qp�ʙ%���[/<��]V��Q�\�$ ���6֙����Ah#1��rP��V��h�j�����k/��w]���Ӓ}��z�>O�8��/��"7)0c5B>�Q�JJx�Y�׆�\{y���J�&���,��M�R�EI��Ky��JNB�.�� �7��>�N�\��#�ݙ�:��M&�� p�:�Ly���Wp�n8���{(����8V�!���'�������=��A4$R{�c�������`yz�TM�F )�,�Q�����D	m�`J�ܨ!����{	Mi9K�J*�l��s�8�&������̐��OVʐA��1~�T~��[� (=Id[��@E��r͸s.G͊��x"e���m��Mi�J��N �߷��0��I�C��L��x!��W�s|��޺��Za8�2g'9W��s,	��ݙ�4��\��3Ok�heDB�4�ġ=�h]qD�t�[�U�`^�oL���<�w+[Ծ�ʰ,�W�i{�`W������Rt�A(q�h���5�Ɇ����"�OzN܄���0>���o�L�c���z�]��n�&��,�G�<:	�+�p����=�m'��H�f3�����#��L��V�>������ь�E�!�3�^Irl�	"��)Ĥ��0*��7շ|�B��M�"ת�]������0X}��24�8�� Hrq�A��2��H}2׉ʤt���i�����Jg9��_��;��D�u*"Dy[�kYIw�rؾ!iSm6=ڿ������jV Q�h&nGQ�$v|� ��A�����Ϙ�g�9c�j�I�E��T+К�a��b�e$�5p,���)g�h�������j' +!�p�縕�T��Anr�8�D���N�
X�-�kio������[�v��<�%};�z��Q2��'��������x�v�L&���^��,)($�)�����'�I^�|��!]ͅ��Q]�岪���^ӭ9Ea�U>O���)��ޒڀ�Z-���>�6ն�8(� ����E����Ȱ���=`�Y�=0�U͆�t[�Ϝ����n��#���� ���MwHﻷ]#@��x_K﭅�;��|��*ˁ,>�F.\b��"LGY ��E�*�Vx��0z�
*v3�z(�\Yϥ��D��y��[�S,��<�%�c�F����1(�4B#�k�Xuպy�C~m�N �s�ǖQ�-K�^���띉;u����yt�% 2RU���0�_�teG�<ў\��bl5�` I��lU�"(��p.��K�#�.���j�{Fv�����(-�N�+������stWK�����b�2����mY�C���M�ǘ�W�Ґ��Κq篚6���� �ٰ�����)Ex�]�~�n�JR� CUF��W@��`"&��˭쎷ԥ�m%�����U���D�@5��]]��r#������>Xk�̀�V��l%FKy��[���1a�p�UiA�����ǭ(iz$}J.�ì�\Pt���!�����f�MZO����ٕ��i�	� *3׸J�Fd�Yjf^��G,.�v��f��l'hI��:8�,>�5P����U%�7wa�9`(��`�~����Uq���G�e�j����d�dȹ�'ڐ��t6Ŝ�`�*.�),�v2�wU�P��oT!�9姉#(�<��4���_$0#T {)'������V�N����-�%�QT=��:y	�W��{�G�g�M{"Nxz
�9_ی?��x��H�m��fJW�өeEQ]2G���q���2[��E��9����$9)�G�$Ο9_w��/}׸Jo�+���&+�kB���-ui\g���X5�i'G��N��yiq��ZdW���;�|.�6$S��-�[w�$���|�y[�3�?��q6D�\k�q�ֲ9y�����g泌��̚�8��Z�n-Rc��X)��i3BW���qVx��5���T��'T�([�/�=�V�O#��b����p�䛑�Ϛk��EnZ�u�1P��m7�wT�RX��z���GPg���%>�X��؛���O�hz��޳����Iב�k��ZH�E61��L9T!%�R&�I�z�*[YX+�xL���e��Α?�o��K�_�w.TD����4��y@��dLw
�Scin�un	6)4jh�x���N��!\�jS��st~S�lCk�O�S�@�O���2d;	���iV��z`W�Ӑ��
�NSm$:�9��F�	K.I�E���2j����7!
��w(F�wO�gu���}�H�b������o�����4��U�����qw%��XzC��~`1Zˢ�SJ� Sp����s��K���*�Rc��b��A��K�c���N`��kn'�&wL��`̱�ݑ�p��\p~ڔ�#%Ґ��#5��4�g�B�\��I���� ���9�M���4�z��:~6�y)%�/�'E�#�sS4*�x"	�u���tn��fu�Ό`�}}��I3������I�%�)+]J��p�?�w�Lä�"�V�g��?�_u�Hs�S}_ʸQq����'_d��a�ڙ��M"��ց�RhY#(�����gq�8o��i���[��n]�I�ɯ9�&� w��\Zs{m��r�<`�$ f��4�����K.
�˓3��p;����
���8RcXp����k�T�K���%��*�澅.xK3�s�����IN@cW�҉j#�v
F���K+�s=%�����{�+���ί7t����M:g�6szd B~,iDdz�ZYbq����}��E��)���JFD��{cQ�H��~�?e���S���[7�d�E���sS{�~��6_#�IFc���ԋ��,�5_Q�	���.#|�}f�ߤ��aD���='�����(L�{C�0i�pJ�u蓺�[���U�<�'F ]��$P+@}��� S�|~�����}0�c�ߔ���U@\?���(�f~��C%����om�+ �\�� ��~6��pN����-,VJ8	M��/I���m��^c=޵@��N�&8�m&��%%:�	�$�Pn(����)�a�r���F�ߟ:��{<D/������V~h��F��v>����c_��dfn��Z���X�Դ6u0� g�Ce���=U�r�	6�L�V0���t��~�����R�Kږ�� �rS��78$�.��EwoHO��m��mv��Sec[��q������:;]b�KI�� L$����\d7��x�;�swnN���Q�Z @	�y�E����5��āׄ��]�3��;_�t[���0�E2��xA���a��q��*��3@�ײ��Y��B����.']��`P&��d7)�/c��1��Qo#LO����ā�����҅� �V,Ci��#k�(Q�?Gy�H��b�1�U���D����=��Gʭ�r&��t�2��b���\Fx2�)�m>;\�!g'���Gh@��NB���y��6�3��L�T��ʬ�q_,h�r��՚?�5F	��3�آO���4��0����1��a.�>���H���~���Lx���C�c�r	m3���cl�4˨��=xQ~��<,�,�|�@Z������yoX t� �>�j��\��fQc6D��u:U�����Ș5d,�ܤ���&j��S���ǖ�)܊�@�ꝗ'R�@�Y�J\۳Q�Cw܁��28>
C	؂�3���+RU��pu�s���y�9�������ܚ�	���O5�֋�Q�V��:F��bZ\cQ�H�O���B��V>q���3M����{�]��0�H_zs�Pؾƿk8�&�i�"�J����&K��
���AȂ�]p@�l6���R#7oH��~,�� ��	E�+s���ڮ�-����۠&l�c�����5� � ����W ���hS!���~_6~~�zd��f�'����L�RJ���(=��t�.P�/lC=}ڃ1�8�	g;(�����+I]��¡��t��@�t�pl�-|�����fj�4�s+�*���$�B�9Mr��,$�ꬕq���"}n�t��u���|��
���(s�4�Er)�!>��rU�I���Vpb�͡44��R���d]�Qo���F��qn-fї�\8�m>���I����;d~O�����7�<�)Q^����ҽ]��e��$"#�}�$�bB��y��]���0�"	X\D
�d�"8@�D5yg���q~s���Rc-5r��7�}�v�EB��)��<H� #
�f90�~%��7Y
v�{D�5�mo�;�䦅�s��a�6(1�6_�f����~B�cT��ߧ�G��4nłf��A�UVz�G��HLep�@|aa��Vr-]{����L���^�^!�ڬz������i�{�0�����N�Z+v'oy
�ڛA_�BC���j����T�Ч%��yp���I�t�����6�]Q�4�R���Li���gӓU���:���T�o"��(���.���0|�}�6ʝ�}��?s��K�M)�N{�x��&D��v7�X`���F"�h[�/���]]:��/ �+�T?d���.�R.Qk)U�W��%e$�tAR�:o��T�C�Y��qؐ�@t�=6�*�Q�yI���i��,z�}��!Y�7rEC�0��#�����8)R���������[VA��O�w|+A��=qK��=�z،[�<��n<BUmu,5{�8n{���k��	�;4�V�l�6Y����V��C�Z,��dd5e�R&Q�mP�_1+/t��Oo\Fy����ǈz#��'�5���
����ø���a���/U�֌��6K�h/�A)��[d�9�NF��1I��ΕN�P�UK����md�{�i\k���pF�K�D���=|$+;�T�]3Mo+Y�� Ӂ��(4n3Bv����04[]���n8��F-e���(uH�Zd�\"�Y�4A
�5�U��\�	b`�$/O�����M�.׋���}��[��)-�J(��1�lxT�oqap�@��2����;)"DT=IE�O�Y�a�� uN�=���!VF`X�i"��R��Apڈ3�죽8�Y��-�l��N���m@�T7�꽭]�#|��k��2Ѐ�_�9����Pz��D:�$ν����$ا!k�ih>���
eȭ�8s{��!IhQ�9��p�*6�P7D��FI��A��@=�����=�Mj[�!d��u!���┎��n8QE����L�g*f�_�eJ�`�Y�b�c�X�Z������ 防 K1KT�v��܁d�~^�V��M�B�R��w�ȩB�}�k��w�@��Iw�n�8�2�k��@��a�0q�	P@�9��G�� �F��0{mZV�b o�Z�:����詚5ّ{�o�N�R�{��Ø�-��ñ��c(�I*�o��/A��P���ZH��í�(7��=3wK.��f�
�_����:?�	t󋙿Of�5�������o��r	�p���Z^ЦH^�,f	�T�O���ᰫ�4��. �%27Q�P��|?����k�=��~�;]ڑ̭~��x(����*���d�x����l��F�Y㊖�=f����w����P?D�:{�Xv?�s�����Q���[�F?ip��=h��D'E���q��j�P�H�%��?�u�.f�M��W<��}j�%�&��&�o�2B��wP�"*�:��Q�NW�z�z�~��vG�M��
>ٶ_��*&;"�M�u-V�9�sw񞚒�)<<>[�5o�gC�(t��پ؁*�L����r%5LNN#A�0�SV-&a���I5xuc���꬙��53�-K��G�H��Ɩ�;����9�+)]�i��E��c�c����@���Ks���M=��k�0��e��%$�ٓm�k'����͔��d"���3��0�.�.��u���e�0�\V�G-��$GFy�P�����E;v��2����1l'mXW7�5X���%��t${��6ˑ!a<'����1�aO�1��(BJ�Y<0�5i$!���s:��,"�����+ ;��2x�%����0pw���nn�%e�
v�_��?���)��rQp�d*Xm���6�����+J��#���Z-�_ح>���;�}�ZZ��n�P��0V����j�'���5�`G�>jUj��;�p���	Y�T��q0�ֳ�Oa׀�0|�w=B6��Q�*+����5A�����?�x+�aؼ6�)_l�7p��	��V|��v}t�/��8�n��t�~���><�h�[�6Ԗ�ȈI`f��Ah.����ar�]�!e8wwϚKx�g*ǙpoR"���������Z�T���6��>Pڠ��~�0�q<7�d��
�yΙ��
a�2�� �1���xB�zf_�E�6�����/���K�|��u���gW�~�b��٠U�
(��ـ$ؕ���©�~T���I+��]���W�� �H�6��l����BK�ܟ���W�%[���$���c��^Yn�A	�ς=[h���JT�7towO�+�� <�~�<1�]?�^�S�x���b��tK
h�OLm��(2��Qne�x�y�@��,��"s��z�������B�B,���@��!W}Da��5�҄ߺ*jf}f�����GZ���(�YM�A�I{w��D"���J��.酒�l��^�Lx���Ho<�����Z!09	$v%w���ͩ��B'��k%�Zʎ��!����s=��
u��q��(���Yb�ҡ�]����������鄗��i��1=WF����DXRl��sX1T�h,�7c4�5��Js4�m'6q�DK<mi|����L�Ԡ�h��aU#�^�v~-pT�U��z4�L�����C:�nhk�N��nP����qW7�<�h��DgZMy�&e2��x���I���P��}{�j|5m3��"8F���J��
���V����	}����FW5�fXЦ;�@U� �*��,o@(c�&M�&z�\�J��m����Y[b+!��5*���?A��te&- ��+�?Q'��uA`&�J�=�.3��� I8����3z��m��T-d����.�|lbyZ�E�NP��,�B��,s���7��|�Jz#�ߪG�0���f��o���%�Q��1�kV���e2���ؙ��T��l��evٮn�^.^��I&�F��+�0�1%��'L�N�L��O��D��c��n��+��).VEN�߼'��4jd�P���c�Z����� 7�YR�q�r/��#�c��}�)�THu9�/���@:�h �ڝ�҆����B�u�����X�'�f�ޟ�d��B���^"��z��И�
k��t�������?
���Nf�|�T�G�+'����ǈ�"�
4=U1y��$O����~��?r��8	#����Iۏ�['"����F������q�Z���7���4��p2�.F:�8��u�木Pl_�*ce}�3��[J��$���4ѩu4��\�� �~k;��V�?F�oX8Bj.�,�����v�-O�r�moL ������s�_�Ё��pW���L>l���/5�8�(R*A��*x_b�Duݾ���_����8�K����l��"~h����!��ݛ�r��=wJ���~���Eʊ5�,4���Ƴ�a��'��Y_��������fy��j�{�3���@՗S[���p|�ɛ	1�eN�6�\ �08��yOw>{G`>�@HJ���� �֢*�-��s3�բ[� 7�'���4�����)	y�E`�4NΓU� �]6%+�5�;C~oE4�BN��jd�q���l�)��zh���/�hh?�^@X�1[�����cj�x8�y[�&(C�@ڋ6��J�d9˷>k ���U�˞^sվjؘ�.	{�D
B�|mq��KT�y	�R)(�X8
�"���N��|k)p�j����$d��O�BW�K��{x�9yі��?����r|v��kR��	)���Z�ݻv4>�F���EƗ��}X�q�������t��1$.�ɚ��Dxwt�I�W��VV�$��Q��~��+%��+�L��Bc�QZS������6@4���\w爱�+fX�p�\nD�a��,n����C�K���_/�\��?������9^}�Q{�}P}����s�_��R�꘲�����jw�$��, �̛I.��:Zp �v����˱6b8ꓳ����.D��@��m�J�b�e��=���&�+�Us�����w�Vu;GDNK�Zf;��bGy{�tuE{i�(����C�8���G�pb�yOV��n��e�(e���n��<���>��m���� �_9E�Hv�����{�@ �t��c�G`�V�p��d�0]�����T�?fI���+�jp�'�5�j�_��U~' ���S9~HZ��?�Q�s��_��=����ۄ��)�����Sr�0"�;Ӭ�L����J��+$(�.@�"8�΀$pN��k�!��!�B��F���e5��&��DL)R0�'p���QT�m/�ߺA��t�Yg��Bl�+?p�n�F
�HTۼ�Ü+�5.�YNBO�`�>j'��A0�_�EZ|[��ati6#���F�)�A�l��������%��H��䞬���t�0l�#u��lfhD�Me�\D��RF�7Q�F!��j��`�ym.qQr�o�V��X�"u�:�X�1�e�n1�"I32 |�M��}���O�g�Fszy{�V	lA�8Bؘ�n�D\�#��9�WӢV��77�`0�A���}��#`{���&0iN΂ 	�#��6$��P܆A�C-<䬃M�Z����E�k k>�K�p7fd����7�3�sx�9�����T:�蔌|;Ǟ�ڮM9�_�y>;�뿋�k&��}*������6{f�;��#�,tN:���Mm�'t���{Ŕ{�;���n���􀣎2���/H�#��@���nXq�l���p�y6�f?�4�|$��n>��v7(��-ý����3ʪ�og��R_�օ�&�%mX\c]��Z����G�=���p�͠�8� 3����6廊m$�y�<�s�Iw��lI��9h��9z���RZ$e����{b#�Q��Xz;�Ү��y���5�0����+���'���H7��)m��|Ɩu��K�*�ޔ-�}>7}a�Bn�&6�Fh[J��t+Ӏ��X����V�<�@���]��;c�9Qȏ,�Ix��mD
����k��K��>���w���^ڰcs��S�=�+�7�����Q��Q�*�Q?qͥ���~ ��6m�:�0�֜�eF�	��0	�F�c�7%�Ļ��:�Ɋ��)PLS��x��{�'f��Ta��4��T��7`���(����Q����FA��_�T��)2}�Ռ�^'�{����My����*
�¤�]��#�6a�C����貞"_���X�FA��9,j��?����D�)�N�%ά1w<��#%ޮ%x���2��d��7����2�z��.#�I��-3rlB��>3&_[D7<���α_�z#����F��r�Ӎ1��������(�����)j.#��eek'j��e��^���rW��oɒ~޵�Kw)�ۜ�I:��S}@���C�0��
t[I���Zòc"�J/Ę�4zae1�g���f�p��Zd`���Y�� 7��X�',�񟈥d�ŊH��lCTK>=��P}ۅ��'t9m�B�:	��� ��/#^/��(��YI2���S��|���xU[:�|�J�y^����T1�l�0��u}�
s�ǵ���2���"t6q�q2 �H��of#�C�|9���ږ>xn�{��o:3�󹚚��a�46Cn}�Su�f��J��b}��O�+B��D7"RqL���Taa��eaʓ����o=��|X�s�y�v��������ԯf��h,���	8�͍o�M8��_��bdjvH�G=�u�Ѣ��:3�E��N"��M1�<��s��"�piVp���6��}e���K~�0.�)X*J�V��p��Q�dT��4�b�.�"��﫨z�c��z�KaHYAOQ/(�wԢ}_�M �ɞȚ����_�+"�$�:$�S��iGvu�>����Ë�k��X���bX����/�,�4���E�1)�6?�Թ�"&^~q��� ���4��XvU(^E�t�7Ҩ�m,���J�|�?|�I4b�޾�d�9AU�@�T����m�����w����c8Lg/��RM��3g�w�w��8�Ŏ��#?�~�D/�FZ��j�w��.�r������ڥ}{��y�N��w��y��)�<��av��ܚ�O���R�Ж�w]��s�"ϔ�u�Ϗ.��Ck=M�r������G'��A9�֭\����?Er�k��qx��M��$9���[1.�6��	w���8�ڨ�n��BT��y�3 �/��j�w\\5L��qa��� �z��Xֶ0CZ����1�3����ji(�:��A��x�y��nP��]a���C-"�7N�@��;��Nׇ<�����J�6f!-�2#:����{o��FZ�O�H*���X�b~���^���w4%�`�y��K���vn�诚\�e\�IE��E2$ZĲ?Y��~�Ҟ����9�S���ղ2D�h^mM�>|�!�
-�`B\���h����:E[�X��>2���%r�?]|,��ߟ�1�rq�DO�_�7�6l��!h�ⷢ���^�iQL���G�G���w�""f��AW{����`�0������制R��X�x�+����B=)���38�{�.�P�m�3.�����u��zZZ�,T��/o�����jf�������r�X�Qb����,/ F(�1�HX1+L��8އ�[ ��C��>EY�w3{��|��A��7�����˖l�� ���`��u�go�$�b�]5Rf�m�ӷ����ލ����]��3O~Z	{��bG���A*���R�;��}�X1��f��t�H����/�͠YM����Y�����P����5R���Y�+_u4::	���{�d:��}�H�|���ÃD�KTu<700틻�MK���t��1�{U\Xg�'I�n� 0P��3���3\"F���%���0T�k�>� x�<7�Q��3�"�\2���M�K��i>w���KrƑ$#�!��"�m]Z�T�%>�f������a�_������i����re�m#��l퀼f��A�
��]�l��b�:H<y�r ��{<!��z7�����W�W���Cl�n�55�5NdK�;����'��` 1Q�D����b"Y��<�Uh���O#����;�ὰ��� ��p{ۑ��_��qe��C!ʸLQ��m�!8w�]�y��?��,$�rhO���^�sՍ!��	;���CL(��3�~a���<G�_PG�z�Fn_>�s��s؇[��-�1�ey��/��U��u��A~�G��� a��e�1q�8�"."��4m���CM����s���r%�/��F)2�Ԇ��s��}�����桬7�j��v`IJb��U�)��
�bo���%�%��a���[��Vq�N}��_�H#@O-�"�����!ve�f�O�T�(>Ψ+$ pۿ%N}�
�ߨ�Y��;�qZ���hiK�����&
��'�,07*m)���N�X��C��r����h�M�yۄ�~��Da��Q���;{ɰw��BڮwȠt,�36�܉s{y��8hy�ҵwg�ܲ�~�{@U������4 �H[ؿ���H2�
�;p��}B���z/�{~�Zr�-\�~L��$
�Y���4��J�r8�������W����U)7rpM�x�6����*�W����Da ?������C��q-�'�fn�C%,�������$}�}��[�����,oԪ��j�Qd��r:�+;%0���$]-���=�鿵h����	/%��u�!��}oS�$�Bs�sf2��֢��6���,s%뛃}���#ũG�)��0���ѹU2���/x<ک2}�}��J��IR)��4��n�FH��CͅxR��1�����~�ϋ�t��.~[T�,���"$K�si��N� "O�@�0~� 9�F�������Oz!�Ad��u�4������T���H�L ����"����n�O��������>[��2C
�C|ޤ"��'LѾ���i�{fi����a��z��ރLs�-Y:�fA[�>�|=�[<���l���Z[F�{�,�j���<�. oҏ�H[p�QZŷ���3,���(�P����$�],��]d�_�����������/ؒ`�Fd�V���JfP�_m�]�g.W��l�KS�p�:�%�-�-�:U2�`���a�d�ŵ-s9��tl���\��L����n��~�Z���)a="c߅�]��%����Ӑ�s"�"P)��5���\�:�[�:4�I�Gp�]��Yj�`突f��+�EEèJbF���f"�{a�V$�ɑ�	��oS|�g �H���'��>�V�>3]��g�J(�bg����f��^V\�0@�����G��%\�n@<��	��K�C�v �'��4��A�fa�Ba���XXlxVHYEB    328d     d30ǶaL�����_ڕ���<��*Oo�?(�%�[B��ŷ���h+�g�d�+�{�}Z����<�����,I���Mjn0�V�JɄ���3�:T��a�yvH/�Uj�$�d��6v(]�,��I]��fA���T��P�Xg�:���b�:�	�z���"��|�C).m�4���h�j�pJ._.�p#�����Cd�~	��=4Z7��4mBT�o3egjf�ul )�#����Y~� �����K�c!yP�P��_�w�����I��a�s,���`M e�_�g��k}BS�I�����j䈇��Bƞ�m�����4�4�5Gۧ����v����Pko�bCg�����t�����x�
SnG�D=g����&;i� ���uIE�������V�����'D�m�`$��ەN����w儆��(�Z���K��� ��-9��.�5Nd�ϜF�
�,��e/��	�W	���h�-:�?�j3eɠ���w���3bZlc�������Lk\U)B{R>�(���r�T�>[���ګ�ߧI$�}"Ҥա'w?z�"@	�F��%���@e{���D^	��.-�_1Y8ɂ���M�����fL��@��M�V_�P�Wn���:�Y�-<�&A��:�K�̸��K���ݭ0���
����3���I\��/#RtdМAр�.���]w�vIU&t���!�E�� �EC�`�W�#��w�ޓ1:��w�@[45B�,3�����H�=ch��{���ؐM��R���R O���sesem��;5{�H|�*�ĳ���؝�EV�
?��5����D3���!���>^Dm�3-�){{������Aꇇ�5��[�;��>%9���3M��!o��Cnx�x������a�j4Ç%�8��E(L��'�kh�%���3���/hV����"��)ξ�9�.��n��W��!�:����am�Y��?�#M�_{<����v��7C��~=БFe�$�>j��$�i4��`�9�ʄ+��V�Q�,�:�)�c�S^�T�t�Qz���#�dU�xy��"\���F��j�Y8����㫎���0�"8�.h���@W(����b愸2�R��)f��f��5�X�Ŕ��RTs+t ����k�͌��N,A�|�X��J����D`����sk�UC���-b�|�dM��'/����\ ���12t���G�Gq↼^(�ȵ<Qj�U���g��;B̝�gR�?}DZ	O+qJf�}5#!�\Y�����;�B��>�ڎ(N699[����M�	������]�X������\��ŧXL����=�U�"��ÿLs�Ll+`Ԡ�`�D�ޭ�X�s���u�oG{�[iE�$�vND�&�ќ��&R�%�C�^����2'i3K�[��Ua��3�PO������$8�%e���ˑ�׍9(40�7��_|�<�����Ԗ�w�c��1~���xO��1W�Q�e/�Dk�-�����\n4*F��B	+;9�9;�/|t�1�z��u�\�#��G^v��+~�Ź�����+m���q�a�`q�ȏ�4��&2�} �P�Q�ut^�zT�U	qm�A�1{��S���/ %��~H�z|kS�u��N?�O���[o%s����k�����Q{�̘z�{��;�\qtD��o�@��b+�U&��I�|�����z�e�^��1t?�$zA3�v5f�c�f^j��~�NX�tB����Z������y$�S� ?�<������2�wa�m�����#��dE;�����;j��T�&�6�ތ�DL�t9u��3��0l*C
�՟. � O�����$?
���>@���C�����#��(c�|��`8"�p�,�I'�Z��7K�M��(�+�WJ���8�h+��QJ�4�` �W%��5��*�/�~��F�U�<1|�eB��Μ���o+l�M*�m]�����k��R�ߒҗ� a�{k���Z<�,q ����U�T�rS���ьث�	&lZwsK=��]	4������I{2`H"�}z'�xK��(�.bW^�J�-���n�B��?��΢s��Dny��[��`�J��oǳ)��Q�C��<�:��]}߾����x:�X3���1�����`* �b�ɤvV'��]C���P�~��c=�1�h�X��Ȟ3���4ҷj�~�ah�9#��S�H�r|(p)35��e����Q����W�D��\@Ī+p�Fy���]�qd/JVy	KZ��ʣ���odNu"ab��������_0�s�O�#�>#�v��i��!��i �Z�:��Э/��&5�qp����Vll?�������[� �`*����$��{$y���<�/������D�e.+ڳARq�����GO/t� _�R:��'[��՛8l�.⿡���ɭZ�g��VC�5�D����p�c����OG�f*TTRP&$��J%����U�s����dyȠ����i-��@K�b�-��Wf�n�o���j0��Jg����Q�Z�1}c򉜏�M?z����ڌT�2���63��O�i��D����j���^��d)c�r���24;A�A�j���;��'#���AH��%�X]f<J���>��pL&w43���Έo3�2�[KЬr��ukY�!��@��G��#\�g3ۄ��l�nԮ�P��Xg?�����^6���y����6r�rd�bR&1f����ô}γe��j���ճ��0��K���)h���E�x�U�R]xC�њJ�G�9�G1g����ǘ��;�]]���J�DS�myq��R�/y����(�k�������4���
=IU�X��>�T˧�7-��_�LF�Ɠ��`�,�I�1<r�av�Ln`��A�|�o�9��9g��(Wгԏ��U��x�$�qT%i��,�������af	���<���$��F�Fr�@�G�M���<U��{e�փ�?Hx�n-M6�a��;v��vI|��I����}��P����7�A�(��Z���ǔ(DA�iﳆ�Ġ�{4�:�*켔��Ѳ#{ڷ{PK�
w� ��i[��X�Y��-z$���c_�8i��ύ\b�CN���C�X9��pl�
!��q!1���kǌ1wku�������I�2b.�h��2���(^�ڀK��<��u�|����!+?^\�$|��2�8��B�	�+���Ѱ�ѝ}}~f�%�}RŴTB|H{���sJp�С���iԭ���S��P�P֙o��@�4=��\T�S���f�8}q,��dM2��5s<���Y K/|TG�Zg��縛���_�@-8}���铚