XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�ʁ����	�~�p�x:.+�Jψ�e����w��(~�#��H^"�$�I�����<��iKwb�'+�������s��2&��2t̻�S\��c��4u\��\.iX��G��`^��[e�|��KC�q^�׻����V���	:��U�+��F#N��eh&��TN�ZP�R�������}֮Z�ʊ�9�z����{C*hr���0G�N��!~2�֐olze( meG���w���W�d9�n�f���!�Qw�u^�^��^$@������/��/U�ws�!?�_ <'�n�!��*�1��	c��^�ͥ���ń\�T��L�6�����=e ,�j���� �A�S�(;k`����Ϻj�յ.7����S�v�*�i�����@�q�n쌥>ê+����9�f�;�rZu�o�����}�����E4��0./�ϐ�.������d#�����YЄy�]�=~L=��=/�Y��k��tצ�@�d��)�� �)3Ekp=o�V���w'礚�>G#cl����%�u��7�\�)�&.	,:"�UI�5�߷�&h{��$��
%�D�t��Mb!7d������۞�|z~05p��н6�[�UZ�,ދI����n��nǨ�*>�ul����,���g�5YoI�z����d�v�;���k��t�l��K�H<|�Q��F�$��m�ַg"��G��3��(b�#�@"�o�"�<�qz�Or�>��̒B$���f>�E��wCXlxVHYEB    1835     9206G����Cύ�<�;�(˅3Ԑ#H-��"�	�MAX������um��N��?VZf1�1���u������NA� U,5Ug��P"d@�����a�ph�Xn��<�Z޷���n�#;�nN|'��\zI�n�W4k-��˙��L�3*:��b�3�@Y�<�E�+�@��3�jK/(��. ��+3�Ų�ˡ�`r�T�{�>R9���e&?�f"X���)^DA����ؚ�s��,J���
3���Cn�|��ޭ���-̀�X�2s�	XO`�A*,	�<���� �� ��ԻE&�'��1$:s�7M����%�U��N�A5���?=��&|�)�K��IF��"����9K���]#&N���4�pDp,��Y'()-����pv]��K����W�;���,E��fM'(���������2�)�~���M��%OD�aA�V��y��|���=c4v�F���K½3�.���z>G_���A�t`�E�~*��srQ�]$쳑�|M»�6��]�\!gI���r���6����Fy�����u�{���7U-=��(DV^s�:.�8!{<��r(�Uy�b�����[�}k����^�}��"�à~�ڻ�������Pc|�o���5������`�����V�����j�)Z�gΔ��M���d1u(��g^9�w�'l��А�޷�fN
.|�e矀y���u��XL��Y"��g�M-��R9�\DJmlr�<2��b�ےK߯���v*Ԥ�G[����� �8p�ޱ���Ύ�pLR�(k�((	��X�58Ay����o���	8����I�D���m��
��d�}E%=�sJ�xNb��l�nt�%;�b�P��C��'�2�.f��?<�����'�<g��P_i���A�"�y�F��~d�~���t1�r@	���Ӯ�W�Y�c���z����\�\?S�ւM��7��i�<�HX�쵣�v�=����_�x,s�����p�F.u�`[Wj9퐀*�@wg9j:tk06�o��Q�-�=2��k���wǥ�z�� �6y±A��i���7ѡ-��C��2�/�g�̮�k�U�����0c��BYѱȕ\�!
�+�$%�L&�VaP�9:#� �_��圏��g�K
��#n,/���040Xx�U����}��I�2: eZ]f-ڰ��S���弎��OcL��u6�B�T
D�^ғX����`%E��\�\}ָ�}����s2z�[\�r��<��FH'��.�3�i%�;�J�̡*����}g�0Y�% C���Œ�8~����k�|a}��er"Y𝽚���EB��w����ek������]�Ol�E�<>��U1��r-���N'u�r��^Ӌ�慺͓���#���+}Rtv�}�����gu	$�Qc��E^Tk�p��
J�!��,%�m{;s!���a��p8�#J=X����|�X����h�/ɡ�N���F�����M��<�nC��[��m^~�G��F䢟R7Հ��`l�{��~���N�9�:�X�o��VI:L�ϒ�;ׅ�ǀ� �yt�Ҹ��K��j1���_CU�&�I��
AP�.ż����g1�yu�QgU������N!��j2ϔ��1kgJי��Ɓ���Z���K_�N����;��x$��J�\s��% #����f:y������;_JH��И�r��:JNq�D+X���ķ�t�B��1g{03�eW!�w��{��@
�|�2j�6֑�L���(N�{��<~�xd��v��&��/o���$8��9��p��rd�S&�G�{�US�i�!��MS�%n`y�;�%~�2�H�Ff���n-���}��u��R�8��w�g�t�k�%4B�O�)�x��TPs`Ef�sI7��/���4L��=8ƕ/�ȡ� �����.x�B�*	0
9t��ޒf�|�N��!EK�u�K����2Y�fXU��pʅ�[�|�{~B_x@kt����n�Uȏ�B�JS�L�-�j�E`���K�@J\�j' 3��[�����b������c��-��?P6�4�ܚ��=������I�_#�^���y�L'$��v��_��*�i:�f_M��3�.J{lwRz=v/� a 9g!Q�&���JP�>���F�1�N�]n�� ���zйnxJ�S&��4�Ņ錎��ꬣK�F�5��Q�ĵT/R��l�c-�υ�_	[�e7�/(�6R����w��Z?����	�/ ��p�c}�[6��J�*����3�?��C�^l��b``"�ً��h�t2��=�d'���,��%�W�Fd.7�X�gzE`(