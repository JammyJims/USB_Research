XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�D������BF=�=4P�6�j}n�J��|I�ȳ��bZ��(�kJt�[p]���̛	+L�§Z��9��Yt�(����n=A��[�{\�?�)�:)\ŏ���,���RV��t����td��C�.c�願N��>3���,O�D��3irݽT��Ĵd3:"7�x})d��l�Lfxt�sffO�B韷�f��S����;a֫z�#L"��Y%|����(c/b�-�8]�g����WNh/���\�h�O���m�qs�Ҭ	�4�@)��*'��u^y�ԙ��{�D�a�#	$�+j	s�R�7�6[����E��Ϻ��KŒ���x�o������=q��,��#�ѣ�y�J�e�T��Fl3��Ӟ���Z�N�S�tqj���y؀c���X�ߦ�8n�����/`\�`o
&��!��լ�3%��_ݼ[!�BY��n�4����W�����p�P�氵Y�i���~p���ZM�LA�4c�e��<n�r��,eg���bUxt�/���pq5Y1�������L*w��aOk
���nT� ~�I�K�v5����k���͆}�t���_���SOJ`L��P=�,ln ܲ7O��9˅ˡ/�b���#C<��ۭ' �A/+�<��;���K(�� w�1�{�f���y��30��Ċ�H�mK�5��)����!��v�qZ�L��)��ViU��,ȏ)��ǧٕ*��|���"dj�k`���j�=�Vի�|��XlxVHYEB    d169    2ad0+M��;o�5�8<������-}nkx��E�]Z�8ͼ��q���Y�H�4)�gՒ���?�c5� a�D�B�^�G���dj����n��VY_�� `·�U�M����~j��)l��z��OYѴ�*��.k����4��J�0$ķ. ޼*�l2��g�V��l�R�l_v�iF� `7U�� ��fl4Æ�"�}M�)G<�	a�����d���H�8�Y؇�&Q���n�����@|��$�'���cx���i]�����p��s�YR2 V�͎u��@mˋ�'�ֻ1�wD_�;�Kk����8�/�T���Ϧv��� ���DN=6���ʺ+�x /S��↏`���v��N
��#�߄�P08�cN�kַ�%������e9�<��z��.��k&������zޅ�+"�X0B�^�F���u���U*�ΞO���b��́}�7���eS���a�C�Y۷qV9����у�o�&��j$���U��E
K�c|�� ���(X�pJL�*�L�FQ�n�S#��W�M��c"�qB��9���$�$
�&����%BC������B�)��ov�,v�x*���
w6��w^x��e�ԛe]@���o��.q��+M^�]T��2�=l��0�wǄ���v��3NP�0�(kH$ ш�$�p~{H�):IY�U6�3����]S�*���W�g�:bj���ƞ��A����b`<f���+�"f�#�E�JՃ�U(L�����2Q�E�m�<U�D��/�1����L�ϔ�و]O��;��{�$�0C�+���+>�#��l��R^���<�]{�)�~I�!�n�lq!t�����P"��r�bI"�ެ�O���n�<���)�/t���4�G\�6O��9�^�m��IP�G�Q;�G��ǘ����槵��/u�QИ�&�;������@>��La�ƴ�`��+F����Ìf�RSރ����8�T��['G΋�7�Bi������QI��J�z3p�!�������q�2��M��/�^�C�RN���9����Gt�f��O��;;%%]�f��N�+V*��ʖ��������
�n�4�d���EjO5�5_��beA���μ��l��dP\uz�r	}7AZvƙ�6�=��= x��^�M��G�St�0��fД��:O��C9�,!m���g�BE���_���2�#2��Ɲ��#���o l�o��	e�ʵѯ*�����r���^V�
#y		������H} �2���D��2��&��W�x��= ��n�*5�N��W��#o@/�S���6�k��(.z֝�ʥl�*U�vg�bb��U���+�(E���/ͪxq��\�֍j^Ҋ�2�#����ykf��S��YOX�|�Oe�j�N��d�'qŦ:6�P?ٗm�D��=��\I�Vr�M��N��m�^���\�6(�$�Qۙ�K�s��rXz6��eYҋ4�02�%��P�2��������R,3�?�q5���.���rqtA1k�e��$�7̅:�}��7�մ�p��03�B���;��(�;�rɝlf�(�!�l@W6騲=�C�����Ҳ��,:wx�:s����a_�g5�Ѽ�>R]Id���ܑ��dնu:�&�*�q=	R42�y����I�9����yo��So[a�G�6�w}t;�qB"��ߵ�J���KQ��;�����Ź��d�A�(��;لo����(�����o�C�5��[K��H\e���L��ԯ���p����	�	�r�,�k��*�V��Io��5�⎞�^��q�oY�)uX�@�ӵj����;��:7gS�����?��FYf���  �ٝ2������M�x�%)���I��9�4I/w�6 v�ĕ>��VPu��+�Įl=o}}L޴ӏ�V���7j.�{����7X0��h�4�<��:�i�"
.���2W�L��Y����L�t�f=	+G�KǫLW��Mڼ����'�ɖ���O{�$��=�xe�y&]5�OZ�o��Ѫ��X���{t�ZB�̎EK�঻�i �̬�sP�dTF�*=���J��]�o}���S�n���NEC��Ћ=)�g��)�:$T��ʏ��QS��B^eb�ͨ�^���]H�8zʜ-�2���bх���R�E!���j�s�ϸ'�$F���jn^Q�j]��:��Lz�Lw�gs��w$�Z"j��c��P��ϑ;��Ү�2n���Eh%�:�)pI�����u��\��u�L ����qE��S�m�1l��WQ�ل�A�	.����*4,���hy������A�9'\x���e���u_P>]�DO���� ��ա�IM���>��7� ŚLj�����dV<���o~k4�A,	l	쫰Owe��̕7��g�y�l��8��2s0E�_�DpG񄔬x*=CE��� �u�l��5>V�A�#Xڠ��]�%g$�"�Z��.�^\��^�#D���C�P�zI|ۜ���mfݨ�<q�	��6�ۘ�� a�ؠT\0����8����V��ċ��ucp-5N�t��'��!�/2	��ڿ�K�[Э����V^�f{�\�Ŝ��CEܶe�6��P_��x�sjR���f�I����ӱN��Q�c5�_r��Y�y�����A@|�T���4���&��a�d����ΰ��~^��}��c�,�X���wG�B���bhL�G���T8�H�8�H�h3����U򥠺˧��̢��ZVg\�ê�NW���c�&�i*�֞�㝘2�M�P������`^g�Jq�&��M&�~>�4�P�p즢��S�D)$w(D��qw�:���Cͅ2�h�3m#O����U"��<��Wuk�3,���_}�*HX��!ь�Y�/��
�)C��m�z!�=2���~�A(�����	@&�0A�S<���6�gW�|��u]*�z1�n���G�m8WY^�)V�1�x���P��&/7)�
5~e�22�k��;�J���3|�.*l+A�?���]�y����T���`�p�6J�m����\/d�n�j��5IY���r�9:|܀ɣt��Vk�����z��r�T20�2���c��1k�+�&?����(Ë\V�������x���Z�		0Z�<��beGI-�tie	�̶���UV�%p���>�KU��m�G&�П�D�dB�SWO�X�g�j=��!b2�1��SM����I3��=	�"uE�w �ԥ�d^l|5��l�J�>Ⱦ���X�WQ��xJZp��x�0בּB�t���7-�/��XA1eLj�h�?��&r(�,}M���NFƗޑQ������С�o��$�H��8�$��H��υ�գL^^���]��Me��D�|������	�v��ƶz�b�v�� L��`+A�B�����(t�_Q�;��������`��-0O�V�v��ʯ��
k�������Dن��F��䡿�ڗ��f�ty}�O����^^F�Ǥg�L��-#O�ܠ�{�y����-h���ԃ�q��½�ߙ�ۑ]�+F4ښd&�3�&����F��<#R����@,y��6�W1�&֒{��	o��H��zo,���@;=�4��N�Ԛ��2Ƣ���kvQ'c�T̵Tn����־>�͝X�Z��	��&���M��,��C2;�xj���p��J^?�R�&����8lQ�Z����F> �ˍ���8�5^����^�������n���?��[n$����'AS��p�F+��|'����Ȭ�jPaX�Vo���]s-DA]�,g*�lʊ=lF����B{9T�n�����8WA7�@0Y�?�;��9^��K~�w�l ���kke�"�Q�;�1�sw��I8iM�y�S}ع�t2 ��^K��ҋP��Q��U�F���RϏY�+���Mݝw��QXYd;�
���YAZI�\B�r�+ŋ{Ǒd��0\v�I4~�|�CC��}����?�/ed��P���9"��z�IA�n������a+�--[���lC�b4nh_�D�8���k|v4�~�nM��ۻ��d�I�P-��چbR�#_������6\J�A3|�Rf��2%��D?̰L�ҳM.��|�6?��@ [����g!q�l��~_��g��s-3��`#���k"�������TĔu�i��o6���D� 9T3��=���=���:�`�VJ�\����Qy�+����f��*�$z~���A�Q�h͐��=]�]����VU��x��;�^�$���x�W� ��)�����gD��==�c!�x�
�{{�K(:�D ʻYӮ�{���FAlX��I�kj��wh"��U"M&�&����×��u�%H�;ӝH�]�jE�*�E,�8��AzY_�*(3���f8�����d.؆5�g5S<� 8�+�;�b�c�`��lZ��B�Nl��Us��;nwxɌ0�����ga�7�-,b�Y<��)��2d�;�-�X٭&��m4�=0o���1mǀ��8-Q�^�r��Su�6]�S�4hs\Dc0��kw��N��Z���ôhp�&i�^lJ���F�{w4�x�&Jrtca�����I���r�F�R/IGrt1�_ڢ�˃�0o[tgk��y4pf�|��ꊂ/��8��xH������)¸I������;]~l�q��J�3���b�V��+K��R�gy��^@EM�_d���fYg�̋��b���Zw����2C��{%RթXwO���lb���6����}���u�?�Y��kN�c���dr��L%�5OΎ3{�So�g�pWl�1�mߟ����D5�ͨ�k�+w�J��ZmWy|�R�E�+u��9�� 0)c�̲����|�%Ť�Tne�f��$auѠ鶻(�j�����IU��v�g�����	#6���7"Y$~���J��F���#��p�0�7�2QAxl.�����u&���/�u7<	����V ]�$[�p�\^�/�
jy�R���h�H~?��.�A�� ��`Q<��>{N����R��Od4Ғ��X�a9��� ��^.HC�"�	#�V�Iǁ��9BD����b�y�U0���ݨ�Yvc]�7�����1 ⿲�*��v/y!�q�Vs��|(E�����a�O�l.ӷQ,�1R���l��Ⱥ�;(��Q#W��8:at�8���?���6s�^R5H?fgʿ�(p��3��)N	3)��B�'�Qb^Z����=(���qu<�)MY'��jkdL�@��3'A���Ă�kŗ*�N�h�k��W�MU�wg4d�G5a-*`�7�!w�!(>���=��p1���faJ�$��A]�E����xQ�����pý�����s�O��IT;�+�6��v�E{�f���ͬ�d�n�PiX�w4��i��X�C�ܖ�y�y�Q�>O0X�_iqr!a�>��Ѽ�����Rğ.�q֐��yƽ�HG�7�0X�Z����t�þ�|�@�L�m�����E,���<#2t�>egѼ4\��nd��a0���]"�r毃�eS��K
z�Yn~,s�l�;�xT��I��,�:�oI��p�'�*���0�)R,[ޘ����:�{����޸����)QT�������r����6�˜뒚Ѵc����E�4�j�(�J��2�4��=�sa�|>���׹h?)B#Qʘ�<a����r�fv�/_�hk�uT�|H��-�TM$���4��=T��OQ&���r��X��2�>�7��H�w�O��KM������w;�Y��SH�0Z�%/it���a)�ME��tχ~<[��Fgjޛ[�cЎ��p�e��#ϵm��⾶H�v	_$�>��	Ɲg��/\&�2B��ի���y�TR#��2_ff�K$��E׳���W�T��/]Ťlgh��W��5��mG]�ӗ��Z��U��|���B��C�N��hWacG=?4��΂�@�Ƕ|��BJjZ7;0����'#�a�ү�k<�(����"��v�Ѭ�b\�K^�o�vy���m�>~�[�F����>A^���)�,���'΄����O�CL��v��~n+�W����9t�2S	�s���-��"Q�>�Y+ݔ�C��(��T>�-�����I>QA�c���L�{��K>+��a�}�Jk�Xz�>Ɛ� 5����rE��48��_W�ຂ�~2�H�Ç2����X}m���qp���&�bV�c� 9���
��#h`/�kJG� �<�h,^|10�ڨ���HY�t.%e�\�����	�5P���*���=�ME�<PKp8s�p��d�.�٘�h�Y��]bp���g(�&�CyB�Lǥx~���d��ۘJ�Y��H4Gͺex��z��N끼�����oR�Ѱq�DCA��)����s�qt��� �g��E|s�d�`�>u*^/Y�NM��+�'ӈ* ~�(�Řh��]�����}v��."�
1Z��~�V�)Jِn��Cc��U\�%�g~t��)PcL�`B�`�/�E�O�$wS?����;>Nז=�����EVj�8'X�W�������gk������7Y|���@��^5�t��ks�ٗ`U՚6��)ai殐آ��V"m�(�rn�1�U����W�(���
�z���C����ȳ��k����|�;_˛����צr-��r���^�	�\����ϩ_-���
��W�-����T"��W�ъ��PH(}Ԯ0DP�i�r���&�#n�s �k���}u�J�be��6ձ����A�w���1P��ڇ��G�;lºٽ���s������I��i�����G��6�E��c��Vi׵c�R�D8NKTO,g06Pk�
#�֘�z1���aw?��Jk�[)�jt��,*�����4��.��Ę����+b��9/�I-����y+U$i ^�A���kT)�~���?jm;�T�C	����@�S��{)�!ؿn,�>藂}�x04^�(>U
)!ר\V���*��%j"�a3.C��WvI2-���]J��	�U�!^��vl�9Y��z��+�e�U��T��;�n�V���[z����	���hÌ=��;�������C�P��ē��ӛy�s(��z8W����GA�x'�c�p����P����v���zvY[A���AcL$�4l�^�>�̓�RUW��j���)k�kI��3���w�������/����+��t�MnC~��y, �;���2���N���[ea^ ���	�<�#gK,l��ŀ�A0}`��@�O����]�a��5A��� E*k\*҆T9!���Λ��O��N~��1�B倧���?�O�'xW��hyrBt1̾�e�*2��?�LH (�������e���G����|4�!�o�"�j�~/�9қS��j�'�i���m�0�lR4���}�M����c������>،�B�f��-�Y�K�ʷ>�����H�k�D���5��֠p$��a|��n� ��U-�\
�Ã����R�ΞC��ڸ��ߜ��P��I1�i6��舟��N65��%IA��Z�g�CoY��n~}I�./���I��{c�v~��w6��e��j��;�/�G6�)�gm\��5��yi��RW�N �3Q��ٟ_���ϥ`^�b�aE�L3ٵ�M���u|q�x��+lb	��H:E��A��~X�޲� ��!��z�d���S�΁{?wɶm[M-y�J�l����U�8���EK�c�Yi����۔�
V�H^�7ޘ�w%�o��K(��|���6:Lg(���
�5.���K����st����ãCɆ�ql��.��f���N���(nT��3�������*�
0x��k�>Y]�D�BG�<G
ř����w'䜓���������j���F���v�_E��wP���h�+,i)����ģV��̾�0f���x$U�w��{/S]W������C��=y|��b�)-$a�V�M;[Q������A��+�'���>�T�-���l0[g���mG2�g���٥����~���ϣIw�4�}�T7l6�J�vZ2�VV{�B��7�<��qy��ђ�fn]�E�^�R@S@�`�:�ߩ���`�����=0l�e&`��ù �G�0������0%%	l;������x4�q�2@6��z���!ѯ�ʰ�j�I��)Cr�iöiRX��dO[�C��Pd�a�T_3�o�'�`f�'ݱ��Fj79�m+�[\���%k����$�*�a۔k@RB=֫��ZۍSv���ޖxT�a�!^���&��B�W�^֩��P�@�e���%e����WT.���T�f�N�26�v���8sb�Ԣ$6�%�ѓl�\{�1�-(N�40	iz �t� X���R�<0�&ᕪl}|�g����hG��ièT���v�M��۹�t���	A���76��*b�m��I��:r�{�wO%^1*�%�G9n
ҽ��@"|��1���a?�IG�(��|k�ސ^^�BTP,��d��"�"�c�HZ^�Ӑ@Ѷ���� ?4}t;�x&0�1���5�,4r$���<�԰��a�h�u1*�	? ��Un!�|�N^ӓ4��-��4Ә_&0>ס�_[Y���(r6�����L�z��8
����)hU3�o_z�M�3����̆'�Rj���l@��0𵱍��T84�)� ��3Y-�ă�Ŗ������N�>>�<��bɯ��#p��7��H����9^�
�ayf�ܳ����#e�&q�=�	,\L��U�덄�bLB�߉�.������oVW���6��o<` ��^���Oc�Wđ�33c�x���]{�3�t�5m	��3N��Lᚷ1���\�r8䍩���O�%�0�y���L�*����"����"I�h+�&5�2'%\�
�|�lud~"�xU����5�J]��s�gs8�-z��-�l�d%�y}�cj�5 ������ѿC�&��պiK��O�������c�-9<�9`I���~�y�&��ë�I4Ir��fX¥����קL-��Y���9\�����9m���D�?��(I+5m�mUp�b���F�g���j+A��	���SD`[�Y�ރC9�)���ܫ1X�X�+��Ű�*��aU�aϞ�I��} ��pm���\�!� �`�/�־v�9k�t��S�)��c�`w�u�g�b�5�����lt�.9����e\bptE�TM+OC�(�WlMY4��
~��6U(E�p��\����s;�TvH�̚�E�x�������|�Q}D����o�^=�ucqv�F%�m'1fx���?�\����_��Nz��?)��}{/����<����㼶���S��Տ1��Eq^͟ǘ�p�+�i$g(^&3t��8���ԩ��Zo9���hJ嗭��"S;iP5������c!R)���,|�l|{H�߂�.��<A��hǝ�n\���ż�Q���e�h����0*
��et >V�bKq����Տ	�w�����.J�6�8��c�!�j���=�j�/pU0N �{t|`��w+�e�9�i��jb*��{Ԩk��hd���c#-HiN�oR�S�"ABEݯ-L��$f�P
"����F:a��.�EJ��G����a�����p췄�lZn���\7x]<��B[��XY��M�����U�;�b_��-_����3n?M@q�`L-�ܑ��ѳQ}�t��A�[�'܊3���k�~�xGC�#��L�̤����o����FU�
OQ�&uN������(­��oǍWm�A�e/diܖG�t��C:ẋ+�eԵ��];�*���Tm�RY���M�ݛ�����������H�}S'�+���X>��$?����-Sb��YQ[f.M�0��/AE j�4��X4��مzV��\4��+�R�:9z�`w����=�5,���卶4�EУ��'��[9�0a���WD=jk�7D��mGf�&�U����|�ĥ�6A6��kLx �2tk!�t�lQ�|��}-�G��=���3���ж�Hd��R:�h��n$���08*x��}��{��llO܎��o7N�k�R�줶�����F�#�T��ꔴ�M����DR
Rg�Q�7ڠxk�z��'�e��{cM�&u�lX���eCV�(��/�� ĵ�
��Gp)�xhy��s�p!F���'����ӹ�w�A2�R`n���̉�)E�S a$��N�e4D�P]��h�lF�;�pg�`i�+�}״�Y|C*'R�
;����b)hЄqa���.�W�q�"l�u��n/���4'�&f\��zs�`\��]OK�|\�	�N)/4J�D��y��]�z�|4���;��)N�^۱��.e�s̃
�{�*|��r�dD>鰟x�0� �e�,1*^��=��O�+�7�ȞWU>�=(���zn�ÄG��j7#��z��sE�p��~���C��A���Ѫ��C7�WL�&�-W�� �M�!A?��Fs�1���)�����|'E��s:$I?�<dC��J���V<#�q���=P�U�U��f?��C�*du�z��rF���s��e����2jkO������	@�%"�x)�M��T%6.#a��~��� �ձS��rXnx�O�Q����U+��t�T�,�hu�Ɩ\fC� |v(E'&|�X�,�?K8'����02�;2�i����7�T�DxK���,��c�#��x���V����F1/� i8��6