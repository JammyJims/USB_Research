XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X99%��ǳ�ȗX9���
,�$^]s��e�X�j�M�"%�YgF���Ȭ��G�U�6���B������[�4����d��T�hy �\^gཝsNRi��<q�А��b���~p/��DU�Mɩd[[�RS��t��G$z)���$NH�+.�������?� ���( �Ǖ^x�h�! �W���X {ގ�B�����?6���� |f���|��� ��KXnU�Y���I]��!�FB���yt]��(�q��|����x�Z��ׇF*����.���r����w��ߺȕ/3�h}��8����V��sD��r;^!�D�x,����y�*'��NNX���:��z��� ������W���yraIl��+�\��E������7�!���Foh�����f.L�Ќa.�!5��8rI+����O�x�/�~I���o�mb|$��}�T2URPgU��t��-�Æ����A����#�ju�,F;vB9PZ���]��J.m���[(�=<<E5q��O�h&��m����@�I�Cx��Sr���Ƚl!����W�e��n�d�ǥ��pO\�pP�x?X�Ф��j�*}�y���ױ��'FflEn���*O(t�Ʊ7�c����^;T��=��_F�t�G�*��?q�<�,������f8����9+�HR���g���8d�|N��K�&Zh����;��)����$SNap�%�]���v�GFù�.�h��J��=���[X}k���XlxVHYEB    3c1e     f10zF�=h��qS�ޥ�k�	3�����+��cj�`U���M�������Ş�q�<YG�g���(�
��L������d�h��B�Ba�6�{�7\��d�yey+�!{�pT��'�����^%Pg�UP#��e]'
Mt��t��өC�n���T9j=:.��u�����MÐJJP��v@O(�G�'�9	�S)��p�\�#eKMe��f�SkB@( X���?*���W��L�@�� O��S���Jfc�%4���p��6���俍+q'm��`	�]#��h7F &q2�dӣ�z�~>eKaPM���t����r���h܋�xZ�����x�xMɁ�U-���#B h��O k�l�0XOc_i6�];���p^�����j��f��S[�����b��L�	> �+i�� �Ǻk4<��u�p��̽���<`�pȠ�١��r%�=/��o���FپeO<��u��pk��Ҁ�YC]����6��H�%q������ш�,;�F�|2�w␊�>6���]N"'�&Ӑ
ߖ��Pi��5�|I$��Ȝͬ�W�M�4]g~�q|殝��vO<��������Ɖ-��;�D�ި�^�SZ�ІmI�����NÓ8q#$�K�L��i.&K�%�{)~��Q�􇬞./�� P4ˮ�*k��� ��-�<r[g9�����w!ӣ{$��`1I�)�K�0�Fhڼ��a�h���m�%���TR��1dK��� i��k��Hw�JVn���q�u��_R�b]�g!w��Ujs��h������pE6f����v�oz�Ki/dT�X��!0`Z[��z�L!͹�@�����2�96.ɻ�4ޏV��6�	�K+����/s7<��pb�oz���wG��+��9g�9�C	��.���Ҥaо �p�X4�b�%:��G�}��=���jI��(��r�LD'#w���U1Z�����t%��Lp�W0�6�;��w~;�X��o]{GZ�Y���v��h����W�%���3E�9$�į{�b���d�ŀC�d?0B��@=uӴB?���wX�Kbd)eX�V��N|~w���>��(��h��ɀ�39�Җ8c�>��	ER.���nH��,�����f��4/�C��>F�N��<���Y�!ɋQͧI�?��Nr���_��Ŝ.c'C`8,y ��d?��L�k�Q�̣-��k�E�Ucզ�\�r��@iҸ-4���,{���c�U��,>�٨�^�H���Q��/�Y�z!?5�Vd�qEX���M"{��C��?�qG9l��9����׏���)j� �{"�0{L���m\�0H9����k�.x�@{���N�����ԌUJ���1X*̯X`v�6�Xm�U�h��f�-��� ��.��-�Pռ6��A͆v���6sJ�ü�3�3��5�� 9��>O�BKBa?��
s.U8�Ie�2�߽Ulֿޒ�k�eP��~���~��.��To�oF�����'oW.����E[����}�:���.7V'�U�(ʹ*����AiTC���zv�-�sҪ�ш>Ƴ��x@���S6I��% N�Q�.;2%~�Ip����d�
�Y����S�A�ps�'�q=on���R
*q��{9�>��a"�Y s$N�A_M 0V�2�	k���CC���^1F!�4o���m1���h��������İڎ���N�6�p��e�����o���sw�˾!�\��9�&�ѕ醭��
�qD=�����W�Đx]�?�G�>���*r(P��@�\�;�H�ʸ��x��\n� mqw6%�o-?mL��TVx�2�V �����Z6-ĭ��}G��_W�q�*}��G��j�"��BS	� .0�C豃c��3�k�,[2]V��ҭ��Q���@� ~�ʶ�:�K��'��Wb�M��Vl�{n��%}�tܪ�������EkVݖS�|H��7(M��wJ�H��A�h&���(�T�*��OEe�y7hl4<^ϫ� u:���k�B�A���zQh�F)�8�����0v�s��pH��b����A�b��w�21�/�W���n����m�Z�Ϟ�\��r>k�_���r��U`@FR.�(�R�@�s`�[�{C޻������u�؈,y�ȫ^h�,M�&2����2p%Pq�*���#�$[�.��/^[1�c�*I|�>+����,'_Ā��e�?��ॡ�4\ؽ��q��,o��8�K���6C��d��L��v���t1�,�U�\�:}R*I�2},��m�{mr]*��Jr����>` �ω��I��WW��32��v��jr>`�H� 86)�k�h�5�'��������h\S�pjp�\�Q����b �[߹r�R�G��y�8X"�T'-T���&��o���e#��ȏPYΆ��)Q{>&�x�����r�~f�di��:���$H9��Q��,����r)5] ��iy��(�5����:Xc�ެX���mġ�q�-긼��]#� `!Z%�+*�n�X=y����@�F��c��R�E��ӭUQh��n]�	[���|dH��д��������L���)o�o2Xx��D�{^p��s̽��:-&�5������Y���Hzô��A*=(�U?u�=6L e<�~Q/}����MY��o*��b��*�pQ�s`����U4�����(��$D~ ��Q�Y�;�h8fY)��������Mh���آ.�es`��T�*j*U4����L�h+�"�ܴ-�'�8~l���J܇��aS�#������fta�qh�wS�i�DԦG�8|$�U�V(n��{PoG��Jѐ���ى�¼���B�E�c��C16��C,��|_�=�:�߅�!Fx�r�il9�&�y!��s�FC�3�;z>�ڑb~Ǘ�<E���*���J�)�p��:Sn~F�ڧ�x	���l��#�a���wd�Ͼd�,U����b=8^fԪ��l�}z���I���0�nF>�醙:�ٔ˨.I#bB09+m����6��+����:s�r�q��:Y����I-E�n�0|��g�6��K����t��>��Q�$E�;�V��B�8O�ލ[��:kr�_/���۸�.r*nZG@�R;*�8�? ��.��D2�B��C ��T�!3C�F�F���'f�K;����?|J?ZV's��'��&d���p����\��3��w��/�u�@&���ңt���F������^������~]Yf�3c>]�o������m�g֏c`��E+,t<�L��1OWk��zE='���p����Z��Ē�EPQ��n�6��q������G[���T��j��%hI�%|�*<ȟ{p1�JtF0t%��]�E��@�H�ܵ ��&K�����&^+D����l�W�L'��_A���#��S������l+�T�`X���b%��&ڰ�oT���{%N�n�#�i��>1��ruP�)�qW�޲���7�.8��CO����v8�Уl�<G(A1�E5j;fj�袒���xU|9�n������Jr^~�����K|(�v8�j�!F��:u�;{dF������)�;�y޸ȯC���<̈́r�w�XX�Ӄe����I ���J+�6j`�eك�����ٺ�lP�d�he\��;���(�	���'��C��q+����i���+��<��po� Y�����"ş\�j�Op�����C'V�6qjj�{=�4���� ����*(HN*
�l��T��w�1�SXev�z¿����