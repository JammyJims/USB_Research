XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���RF����Ԥ*HnH��{�e�Z�)ʣm��m4���q/o�U����m��^�݉�᧽��4I�7e�=@�7�[*�l���;����ǂ���w�s
!�}O�IN
��F��4�l�0R�fh`gd4Z}1�N�!еIbꐲ?N%;��R4��Z�	V���|�:��W�pb2C�3�>R��ݲw�߹l*h�S�!�2y�H��f]M_B_��en�H��h[�ם�.f���jq�fi�|�F�ӌ�L��No\J�ڻ�L"N���ʡ3��K�b�K���"��DA��;���=w�}�[3Sz�#(TMr�Hצckj3M'���z-�w��t���3B���B��u���Y�y�2}����럀4>F`��J�[s�Z|�h������α�^�XTe���u^l��}�s[�bᝀ	���&���I ��YrnW/�(�ō�2���Ȼ�X6䤋
?"|�3� � �N�)��3��.ӌʵ Ü��|��/f��Чt�N�r��	�>J%T=+Ƭ��KHP��J��[��m�i�cr7e+��uR��֦�o�M�h+��:I����^�dq�H��Z��nߜgj́�d�qN�0��τ�L~���hg��q��'ķ�QL�o`	�>�gJE"�1����}v�7E'�d����� `���^K�����{�E{� �#�,��%x�^���SQ@8qH����#l���+X�d[�I]�j��Z����׬�kΙK�IԢI�XlxVHYEB    2b07     de0Q|-KdCZ��AN^iE[A&j5E""��X��s���ȯo�A��!e#πۅ�>��y[��5I�|���oI����]m�p���k���\�����6�A�\�o6�`-�)D�r}��'Q�,댗TZ����)���vkǝ���v"Ny����%pl�I�c�� ���V>A�\��T�� *�:;�%(=u�{��Cu��jf�!��W�;`�����E��������������>�Z�:���)�qQ"�G�ҩH�Ò�TJ��*�J�5�|�:���<=:�g�8J���P	K�����w�s�h�̽�C��eN<�c�.Z�sCu�^"|
���;���P�?�_2�^'�$Xm!b��fG�0N�B�+�	�������H��.�c�(���rrwo�?�=lS�h0��J�@������l�r�Ә(:I5����Q���!�RF�G�s��۹���Y;_U��vqR���PQ��ę퓋��}o��p�x(zp�-w�f�Wf8ߘ�9?β�(��be���}S�&�&��?�t ��v�%^׵*#��ݦn�b��O]�py��;7��v���5�W��`b`���D�j%�V����2q���N�<���Qt�˫�r\�w�4/9C�ڮ2*�j���9��A��kV>���)j>%���0���rӿ�9@upQ6��ϭo�T���m�~�������[�v�[��`T��� �!8�O:]U*2ఄ�8�w`d�~}�i�f����Bk�gu�E|�7���'$M��8t'K�� e7����1�%�<�p��pÛ��\w��U��B�z��	¾��u��yv^�}�J}�zB�j��A�AG����������o��"�����[~nUӈ.��+ixP	rƹOX2(pXY^�H����t*�U��St׵�����3�䣔v�A�}C��p*�ө9�|�y�0�16����^���#ڃ�,	����7Б����=&�%h�0j�=R�ґ�4��'�������LL� ��/Nߞ'Ft���o�ĭ� ~�Fd��cXQ;=�R�"��D]S�xUԠ�=�N��۪��h>�S��J;�{qh�=g]+͔�_#<�'x=\~�˟�j�WQ���Ĝq�]p�h�������=����$��3(��ta��
ʭB	n�Ԋ��Y��ʽG\5�X�hM'
]��TA���k���&U|�1���	��b^�|�Χ�W�!ؙs�k�G	e��_!�a�&�?)g����z�r��b�T���DGxV
l��5��-J�m����R�^%��B£��'�W:�[��_	��D�0'?��[U��h�y[xq�����9a'4xy����2�!���s�
�9Rȅc[�=?�9а�۾��4�q*��:����M�=�f{Y����L��$Yiz{R�)���M-�9�h<'Ѥb|�<nCu�ԄE����9��&`iBS>#q_�_�e�pa�z�H�Do6ׯd�(E��+���E��������l��LMme�&5T���B�~�w4��G�ܣM�Ň3�{�� nmI@��&��X��UuT������!�l��"�H�͑<yڏ��h��`���Z���kƧU��LmYO&K;�1B���#zO�W��De���fdє\�;�)�Z7�S�]0ٌw�Õ�S|���r67�����)n^/�3d⊄�6j���Py����̝��/���߫�--k�Px����L*��>��Zה�7��j}�W��4�m�d(���L*>����>	발�]YN��r���Ӈ>X~h��g���V$5s~���U��c�a��|���S��XŘ����5������G��5���y1| P�	�E^(k9�P�Ma�5�R�fN�A��%�F�v�2\8z,����%Ȋ�nh68^\Z��˫m\�����'��Գ������@�v�Q\n�x�ʁ����S�~e]	q�2ܧ�ˌ�5�7�l!�/�����^��g����`�!��0ޙ��&���������S��[+�=�\�?�Si���  Y���y*��ܖ��\ȑ�g��?_�^e7��+aa��
yɥႵ
'�t�꫊�b �/�U(���8�Q��.�r}��荎r)�|�)'� r�D��BG�sBy`���o���/�8���8�A��'za. s]�$l ���۵ {Z�yk"�1OXz���w})MХ�Z��f�,A�(�g�l<�a�M�AzI�k�.h!8D�����W��6I41��+���$^�Hp)FԊqh��=	��K����i���;.Xې�w�j�6����J-����ȸ+KڰL�p�sJ���]U�2��1P6W�}c/.���|�"�l[~x؞w&a�%&��%� �n�_���VF۶�7��nY�
����*�f��A���n��o���G��p�kHu��0%*/ݖR�gj����L@�Ӟ�<��cc��,��Pf�+�'[�K�G��l�dٗv~�;���9Y����a@�E܉ŧ ����`ԴR-�H�[��i��5�q�n��vp�@�sH3��M��Ht?�t�T��s"��5$���q���n�a:)3�C# ��]�S%>����]b`l�nIݶ��gإEW�$x*�tk��2�$�w?�A���PT/�U_"�9���e� �(�;p�/[�Tg�?����u3Ќ�9��Vʘ�0&U��m��������N՚"g���@��Q|,��P.Z���$�+6>��@��;���E���]g�B�-�9qݮ��Uf"y}�"�ANW=w��!�����/��ˀz)�:dͱz�~�(N�9��#��7Mh��$�ҁY���tZdg��ٓ�l�ʑF�(0������.��g3�t'�\à�d�ht����f��C&�'�����)�I���9*���Uz�àU��c��l���ȞG�v`��y�NCw�`�e��C��'���(+�Fۣ輓�:�D�`Z�N���>\&�1Ze�Ju_��$ɢ��M��@-���<o���m�����B�/�j iM�@����6D��a�"�I�[CH/��b��*�y�T����P6�e�Q��FŰ��/B�i��X6���%z��%R�^D�-�{r���D�ڰ���hj��d����˄d�m
ֲv��X�<��� �KAt=�#�c��'�m�ϩ�ٲZ�=�o{g)T{������Q������Wn�lC�L��ȟI���av�?�y�B}�X�5:��O�ܒ@��������s��HȰޙW9��&����T����C"��Ҷ��T7���o�xdp�� B=nmL]$�1A�57�梲�kN	�r(�#�����S��m�]E��־1Z���p��/���oe��A�5R΍OM7SN%�r��H�K���@�����G4;d;��zx̗����~=����d�jᇢQN�_tW�&�o>8	��