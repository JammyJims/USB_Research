XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�͊$�/��ͰR炯yDlm�_��C-�p���8���K���"*`�_��
�Ì�3Gfđ�,9���{�m�N]���s_����yX#G>�_����e����=z�����:�Z��/��3�+�ٻ��B6RG��nҦ'z�l�^D6����֩�R� ����^�:/b+]�*p��m�ߴ����?�)�ʣW�Xo��{���g,P� ��>M<�W.�S,Ț��j��h��{�q�G�U��,x7�"�.�A�q��A��;xS����/ ]U.��6*��i����b'�Ԙ�n���'v붶�TT��P��"c�.��|ĵ��o��;Aq�ՙ�t�ۺ���n���f�JK�k�Z�W=笳��ԁ$b��з4��N���/��EL�;
�Y{f�w4�zy�I�δ�����_�z�Xft|�S��)�M�I�3LKA�҈�!�f����prk�n�ۜ�I�f�F�,���i}�y�����h����W��p�V-��i^F��vk��R3W�L�\<G#���ȅ_7eʣ�`a�ٶz�*6\q������鼉];5�g�$wH�n�eN�R�5�41\j�&tTHX#�IF�i(g́Krú����j �-��R���u;ɪR$�E\yW�_��y�Wqn�ɖ�G�[)u��G�G	T�S���{$+�f-;'�3��3�v
��o��uw����J����1UǮ�FAgKP��1�x�r�eׇcHk�"��b<O�V�V��xXlxVHYEB    10c2     760�4A��������vTM��힝g2)sCH5�/�$��0���^���{B� K+�P����
 iDZ��w~�j�|�喜?J����:E(I�0�������]�%��+F*�*Q��Qz�:u�"��.OχZ�>��7���ݓH�^�T��[�R��}Y�G��#��w��#S5#ڿ�Q���o�+8�� ���p�q��nz��q���M��F�?
��o�	��:
�&��]]1�p�r�jΦ�6\�`�-l�:��R3��1TH�en��
N	�)�Z��)�W>���,ã���G"���j?�I�� t�H=�T蠫�kC���[J�����Ka� �.��%���.�� H�˻C�2V��1�qj�}?��pl˶|Ŭs}�ʖ�ϟ�u1���<��4d���,2*"�/*?��_�8#PL����i���^�N�J����\�f�%��6�ݷEv��Cx\|4�����pQL
Ö�s'�;e]0I�^̩�%�}2͗�_`��Xw��@�z����Ǔ�9��~�ҭ���NEy���kS��.%�py*��E4� jDN�����KÉͩ�%���.�A&S�w���ɊH�3+g�<���x� ���*���+ݥaӕf��O��q�y�Nt`�ɋ�0ٻ�ˬ� �m�6`y�2��x�fأ�j��;�M8�:%��	f�
�޸��M6x���0���)����g�g�~�ʄ�0z*��Y$�+S�{aJoO���C��}	���3��ۻ�h��D? ��Z=7�픘���V����ٓa�����ʋ����ﴨDUr�nX�"��
r�N����)�uvPF���������-&�)��8�"��M@�<�`����Zr�r���U�Xe�Dl�H%]6.�Imc!��_d1��~��MuN�Kޔ��_��4{�{��[�2P���G*��i�����u[ .��զ��Ϭsc��W��_����YVĠ�V?;�Յ�d������N�u��W������l4�h�󌏌O/x;*�����ěg��x�1�Ě�T�[u���a���2+�Jp.B�F��z�"{���hVW#w��	�!�&����^n�v����ލ����"���x�E(w��O�0�״#���ó|5ɾr�M�w���ْ��ۻ�n8*}_�A�-}��%LZ�\k�.����؍H��3SB�5��(p�����L���'lb������"Co	7�/�s�qñԄ%�ڵ$@	����&�lڮ"ea���HI����:MkLJ�h2ܡRqs��+�ۓ� �$$%=��*ɨ����Nӫ��k�1U�2%��b�b���2���~EV���0)\qU��8���I�&4j�9�|�P��3��������b�
CB�ܢ��+D�7��Wx��%���X��reT��8�tn<���������~�+A��dJ`����h��#!�S�@����P}� ��T������G�S.�S�0�W=#�X"̓_1`���0i�ǊI�T��,�ڨP7���%̢�o$Ҁ �
���*�KX< ^^�=s�,�䲃b!!��Zi����,[om���ʄ�8lD�2;��eW+�$Q�qy���Q�y!��U�_3Iy���2���i�͛p;��Z%%�g�h�G�l�a� :�G������$P���0����V�+C��y1%�ذ�i}���R!1?��=n.\��we���$?r�8���eH���'���t�GJ��[̨�bI���xN�Yj�$���'��!<��<�3N{n�u-�������#�Ǹ�}$ �+l	<��v�=b�
���Iҿ�ѓ!�h�8���Z�Vy�c�X��pG�b^��!�QpOI