XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B8�[���e\���-��y�� B���bI�R�^�.%��ԝ��Ei���Fo�J�b�D�m�)�E��lC	��a?�V���Y�ܮ����!e��[���B@)N�A|��m?�rMPHd%��&����/�6�(m�C�����<��9A�a}!-�Id �����z�����#�1�v�$�I���1����V\�w�>۩��8���a�L��V�������1v[xc���p� �6}T#��!�9ՠ�����x�L�������ڇ7�O���̈��BG'�vE�k�ٝ3�i�3�|���7��USC9�XE��gNޅ`?#sr�"T���k�>|KۑZrFH�J<54G	 ���Wr gs��!6����̀�{i��o��v�Ֆ�ud���x�.��8T(8�����'K��Z��c|�3�4�	H��\� ��"3�B�1.�&:<�Χ:��J��}��KN"��kG~4].l�T�(�M�����]�J�N�l�1'�%������>��_ia����њo�!*�E��q��ĸSv}����C�1`������"��n����UE��r�]�y:n�7u�bW�(��h��%Ҋ/aE��q�e�ȇ6|���N�C�����G+xӊ`J��q��s�p� ���O:}6��O��� ������Ƅ�1è�r��͢�T᮱ϑ���<a��/��C�̋:o`�j��O�/��`F�\�^���~�cQ�_g���r��XlxVHYEB    7d0b    1ac0 �����M�����Z`�C���k�U�_偊.�ot�;RC�s��9kiwV��l�L�����*��=��7��5�񂍶Տ�N�klT���2��*n���F�@���p�H�7�����nA'{|�Z<��- `.��ֈnhi��w�̄����r)+"�s���!��RS1T��wF�zT���ŔF���Z%��Jbu���5ފ.��/<,�EƲ<��.oV}.J^�{�f��T]L��!鸌��dɂ�<J�S3c�K��!�������|�*<�'�X,�AH+�9�;�d�a���q������7��J��?����y��7f��j�x�'��,��%�/(*k� �t� �4��%j���%�a;I����kX<��aio M��A�$ǵ�,	R
~U&k^����:фp1�i<8���l�6���>��ZJu�*�\2�ا	��ٟ�ܘ��#�[
F:��u����N:���9¬�L�6��8#�a���S�tT5���V�M�P������ӂ��	N,�_���Xh�s�x��V�1�N�կ���ѳn],T���{�a��c�n�kh���b�R6�"n�ʵ�$=�#�$ �U�`�iha{��E��I iR�#aR��C�Տp�W"n�Xz�K���AH��M��3�v<���1RO���,�(��Q>�/|
�}	~{��1�^n,�F�������<2��#�츀��-m�GH�0E���/n2�����P�h��� �H����晧�DnP���E�Q}M�A�z����5F`~�P�rk�����5���l�%R��m6�@=�x�G�܃E:����Zdik���f�'bVE&�6Q3�s�-6>р�d�_q���U^L!�)Gr��#/���
�Q
-����X����:���L��Y�֐ā�]�X�F?����t��.?�F�������9aF�ҝ��ȱ��e-Ď�8���-N��NԜ����d"�} �U�ގ"��|Kb�����#������@�C�}|*�5i1�6�"�%�P�w���ZT.�C���?_�<����k���%��K���$.��譙U:\��z�!+��ɖ���=�G�^��wi�W^ d��V���B�%x
?���=����^�6H����t,iQ�ٗ<f�0A��qE�֞�+z*#-�*�E<U�8g�TBiB�j�>/CY(eϟ��iq8��ٿ��6�7���#�!�͊�b�+yW�� {�oڇ.��u�M�b��-���C<�!ʁX��;��S�cG��
�O�g�L�$�D�8d`L��~h: 
mc.{R�������_���td��33r6R����+xB���\n�р�I ��˥:L>u��H������yԳ.�X�d*�����@�j���}�����c�d4P���A���j}���S�j�@�P��e�#k糛����?�g�D.XUG�ѕ������7��4+Q>����LG���8H�0p��F��y;�Q���r�0){q`bV��x��e�����?6�c>�Mh��rQ�Q��à�mդ\S��])�DLFW4�O]��:�i���\��dw/�V���L���+o��!���Cjr ��fL��7MϘ�w�9�jut�T�B;<X�����i	L��	j��:#��A���aL������VtA�'��s�W�)���&�D_,���3�aP��Q�Q��L�_ �xvy8�"�?�6�����oR>|Y������Ki���D��>���"D�a�>����o�佔Yg
K�j���*s���
)S���flBK�_N�wI�����q�d�j	�Ά�h�)2ῷ����(o�wN"�%�:����M Ԃ�ѭ 3�536w�_WP�c����
�L"\��(k4����r�=�/=��<JK�͎�ev}� |izҙ2��n�^�R�wJ�Vj���R~z�������a���>���j|�􈵖��*�{�3�����uKٷ_��2n�*
��� ��BQ�B�)�+��;9�%�Grނ��))�
4��B�T%I%����ٱ$z��;�sص�N�@g�Ru�gK�����z�8��櫢��R!�G�SA�3.z�F�������]]�e�=��hp�� 8�4��-�2�
p����lh�C��z�H����s�.�g�̇��R�XH3c`3ZP�"+w'!�`-��&��%s������H�n~��=;G�Q:��h�<��̣�0B�1����~Q�_B�Y&�h��>�#H��0x�*�
cW���S��0��`��oh��� �b��8!?`��<\������hwY��h��s��^���h�{W�t+�v�#�S�[j"I6-�D�*�����G�*k@�&/�G�Z�_�/����E: ��^v��s��K!��r�FDYR]��/��u�o �������>B}B����Ć.�������ܥ��X�p}��|�����e/4�[�w�QГ,�SO��n0&�l�*�4@E�e�鍙�����L_~��k�y�ݯX��ƦY��V�[F/��gJ��"��w^�����d�)�e|��"��'m)��vو�%�������<Z��l��Һ45����+�(�;���;M�K9Z�pj�bx�ϜS��&��+RL�4`��^��-�����`����P!��}e��y�+aF��w��R�%�ӆ����ʽ����moq�}W6����bٸ����,���5�ʦM�5h���M�d�V��n�R���:ku�~lg�~I5%��e��|�+�|��A^�~�X串vD�
�-�5�VP�^�>R ��?�D��������v�x9#�m$6����ͤK��'�^���q�'�IZʹHC�Q�������|�#���i�"v�6��Z.lǒB�d?w{;�I�\�#������L���ƙ�f/���M^ο�6_���Qdf)��>ns�p�1��s�}BO����������(�d�vS�&�$h��[��`���Ia��������4��\i�{כ�F����K(�x2r�/<%��R��1t��Н?FvQ�a!
�e�͙ala%~u`�PGa�LND��\�S��?�T2�z����5YJ�Ԣ!�C�6gj��r���F��ƀ;�>w>-W6X2g]_�{�$S���iVgG.k\��*�y��Z�&�i`�E���a��fr�"@�!~[>��?F�k]!w�X��5�58���@��ږ�AQ�����,����Zz�@^�?��#Xp�E)a؅��h~�L9^J�?^��M2ة2P8�wF�޶�X9p����*ئ�"��^Ɋ����ӨHT�:�h����\yE?O&bp[@��n�~�X[�T���rw͑�/�V�~5�A��bk�z$F;����̔��E��b��*�k���5.�.��s���Ţ9�I2;�E ���<��G�꒭7sxǭgK
�h��Ћ����S��f�ql�+ uL�P�*��C�A����)6��%f��(������ :Jf�øaH���[�v�i�]�t ް��R��,�/�ׅ��dc����V�P��^�DHu�9�z��(E+D3+�5�p��$?V�R�/D�t��-��1f)yY����L&�=85#��8d�K9�3ie=v��AZ�(�%v4=?>qBV5h�8<A���bC��VS�μϜ��
ڛy��f%1ǹ7�]�QeT������g%�i�?į����"�i@�w�-s�e�I�TE��pMb���i�l�vm��܋�K��'�Y�e2/�R.Q#�ߝ�*��n�`0��Z��RU)yQg��s�b��z�Xr��Y�Y�'Uy¯����+���a�{~rq*�]��C�t���������j-�gR;���4���h`9w�!Bx�A����.�n��#;���Y�����q|�#���8��5v".���<��pҷ�rZ$�W�s�>@e8x��B"��X�B�|�� Z�t|ҕ;C�&0AB@ɿ�h2����[�u3�ܑ�o���/�N�K���N�9̶Җ�vh�������5���a�.��J_�;���V�\IC���"B�A+���#�J��u�]��Y�,�9����tip$��¦����7�3LK�b�ζA�@�ρj:�
 K#ӛ4 �j�:v�e���&8�֒�ٔ��jS&��E��z�^���1'a�H��A7�&�(=@����ۢ��-:�C��!�:��H��%�*�1�I��n#�d,b��WJ��ːB_/��$���=F�sOܝ6V@�
��������+��Њ1�;z@=�6w���t��g���eK� o��h�Cj�yl� =����"q<L}g�t�O��3ې�����iK.�g�"����Ĕ�K�թ688D��� 7G�������`��ќ�u��B�$Pف�B2��>�S�f�I-�I���15�����I��@�O��e�E��ex��'��`	��MѼ0
��-�����ֈ��j���yo��o��Ϩ�l6?�i���P���R�A�s/���R�oה3/Q)=<n�v��	�%�)����+�����Mf;�ƣg/%���\$VG��d�ט׋/�Zb�o�V�P,R��N)�d�u'��̑�%";,�1˃6����(�ؗf�ȧ*���`�ߣƎ�~��f2�u@�9F���_���
A��y�x�. ��'����vk�/-�������~P�#.���=����-�b��Sr�}CD��������M��?s����pd��+�$�(5���=0��b��u�@�Z"�:"&n��ک�e�%s��пŹaV��<CL�������w3�5����Y��n����.]���&�ׂ�GG�7����88���]��{q��_��A<o5��ǍM�˜�͛pS�"P��K9�GEb�#�C��C��E���J�\Ha����(v~�W�VA��<��ؐ�TR�v��`a�θR��S8�X(��1��2s���f7E����;��6����#�*XOt��݅����Ѭ�(B�y+%���?�we�ִw�Pu�B+��;�=���.�C��{���ڇ�n0t�Ȅ�k=h�����e.�����J�7�H�y�)��[CR��z��+vWzb�eX�G)Ǝ H�_��#���Wp�A�h�G�:�"�dG�}�G��JΙ��NCM't5Xދj�{�))�������nFʀ�.Bl�ڑt�[����0��{t`%�w�����3��=�^����ޒ�$aIq9*�c����*��3
:Ȃ�O&�(;��<9t�fR(��HN\~EJ5A��xH�2`|�F8����<QY6q����-�	�P�8��h\�e3!���*\�Ѹ��ᐽ|�����Ĭ&�E�����v�y�)����<Vmй��� �ZP��,��"f>�*��������a߹|6�O���iRK�8��2��4���el9��u2�E���Q��SL����P�/�p���Knh�@�2�?Ny�_��stn���6����XB'��}W(�8-�t'� ]�/m+.���Z/��e�g������xy�e�P�����,�u�3�\5�v�{[�QA9W)�\��";���O8�q엁~4f�u�Q�˲5~�
���<���ԓ*�8n���ky�7��D�V�����R)0���T���J�0&�w+j��+��jݢƁv�t3�к
5gcXU� ���Ŷ��>>����"���&�$�� ���C�����M�Uh���թ��w;7�k�x��އ�zt��`v�]��}�c�i��O���������{�/�N��BHT�hs:�0ꇆ���"�����߀����!Y�=�S#�˚�%|���‴@,MI����[7�L��/�BD�Y���\2��C(^�Wܶ�7�M��)LO�:J�R���S�qg ;W+���?8u%���{q[9�^��Ri�P2�X��n�حݘH�?\7YC6-��>3g��r]�H(<[�'n���?��cϪP���e"1Ƕ��&��r��k��_��w�s�p��l��m魠y�/u]��r�;3x߃Ej��
R	~ՃT�֚,�m���NbwIf��%Ź���n�}�(O�%�5�i�WI('[-���>�V�X<��'$��Q3�0|KtA!�$<���zq�x5��	���ǌG���1�9UI���D��V��8L�]�P��ʟ�''��g=̊�M�(;�2r�����
	Lܦ �b#��Ѡ�����Ǯ��f���z�_�y�G�3�QuPX%�őP	ǆ@@��C8��k+]+I=g�s羙�nCy��k�6	szz�S<v�*��ݱ��%����N;�5����m7H�h}��4�'�RÈ�0�м�hk�k#G�e>wb�����*�1��/������1Ᏹ�������F�/�0�!V+]���F��h�����!�/=���tl���O��zxϪ7���{��v���?{u���e��8��H�f��N��+�|��ZU�^�<�Obr�#r�Z������z���i�T��L1��p>���	`VV�=��;���|3���*[�� j�ō��R�}#G2OH���l��J�7/<4W��%����Q�
��G�oj���f#a̷X<��wp�{ �B�[i�̵.H��]uҴ�O�D��k����Q�����*��Cjm�ǉ9�4�0�����p:�$�5�Bq�#��P���5<d��U�%ȒeEe��w�|NFEݩ�B�