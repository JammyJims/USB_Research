XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[37yA)�5Wo����-�W$kU^l�_��4�;)�ff�b�歑�@q��jk_3�U�4�9�ܛ����mZ/�@(5���h�ǯ�n�n3A�J���=Ŋ��N�6��-�H��2	!A��_rz�d����֧:�9����i�#�S�����%���])���M��G=�����yON��� �ʡ�G����'*Є�U��aY*�����\ P䭟ؙ�L �f��Z�ʳ��6R�qʬ�jf|A&')3y��ج����U��a�����j���&�M���ۯ�/���Pi�
���n�_+oE ������<�'DYȶ�����ɜ�K�X�B���"L&FC&�c�Y/�#L�|��X���b�"�{!Q���61Q'����֑]���܎N�<濘�J�6q�$�AHs���m�jD�9_����z-��h��{"��,�gk��;�:]�^�Hi/Wl��o�䛬���<5��/�>u&y�tb~S�4ǰ��gtQ����b�M�I���42͌�z�v���G�H�u_��h��ř,��z\?��W��3�sk���H�����gk��k�n�Dg�8d��Z��{�\!S8�D��Tz���|4/ɷU�Pmɂ���nR��u�߂(�Ҽ8 �ZֽI�!��A/���3�l9��:����.D�.���ӌ$4�a�ݯ!R=R�0���1py0JWӭO�I�_�z�]�=K�k��-�Pm9aL��[ݘ ⵯ�������B�cQ�� �rc���pXlxVHYEB    24f1     c20��}V�thP�2�?1Ko��'-K?� ��X���k
PZ�#����a.xJ����}�/ן7PN�֖��3�� b�������-�0���#+��g�饪���ub��DU�zxyv"+�}�|[��c�#4T��zI	��ڔ�F~�cA�#ꛍoL0z��=P��ۉ��(�yȋ]T��K�
��(�犙�MS��7�F7Y�crd� �4���h��a�mg��Q�g����o����~dX^���Z�)x�{ �5P����ө�{7\���~��
�zn��Y�b�vɄ����m x�V�r$�yv�:�2y�[R�ն��G�V�����]��w3���Ώ���CU�Uw
	��@�g\ra��a�B�/[Jf�Z��>ʭ)U�������o��������E�A��6�>W�K^M#"ٖ��r��2T9��l��/���%�P]e}��N��m)��%w�ŉl�$�z	�1B��]P����#���<!�nb��'S�#��V�F)�/_N���ؚ�].O� ��$�s�6�aU���&����H�,�R������ϓ��/�e��ώ���&Z���JdU �;�y��Vp�F�@���%��BEjAgzх�{6���=AcT\��$"|Jd'Mg�j�4��,t ��Ӄ���wKƿj<������Y�����K[i0.�􏼒CK�~]
��"�����̸L?�0О�,�2��Wڢu_Y$-�P�6�i�كv���q�t�:)$=�fR���5&��gN�[�au��Qnϓ3`��l�T����W�:�<P��=�O�Y�u�����G�B�>�S�1t�f�#�����K�X���=`7�V-����m!��fb�%��/�cm(pnRh���_��b�,DEM0�e���+[�$?j�.ev�w�Z0���|�Dbj����l�P�ZǊ�A�<��|����ݬh&jhg0A&���aO�s?�s8�A�7$v��y����ra��ϴ ���IB���ա(RSZ�^�Sҍo'���Y·qYz���<#��S��ZGJ����3zfҧ�[ ��=
Uh�tq391[A��c�KvR�,��<��K�#W�b�q�"��uŜ��䳚j��>0Q܇)�X��M������8)�:�=�3��(n����Fe��x�����Y��k�:�����민��G���,O�м�d��En�5�\�s�Vg)�i.�p8KG�������� Zj��R�bD9Z��Df�K1F��\��6�2��+^#�ݴˊz�%�!�떎(�i#�ը�ͮ��R"�f����$��,��k�W&Gk�*?U3k%��熻H���__-�i5}��԰�ǴṮ�t�ފE��SU�p0�^�f��(�&5l<j��=.p=?E��n����e���(���;�%z��g|��c������|ݾ������}�z$���)D�{��������X�B��㙵iU<�h[p�%E��HW��/���۞�ٍl]�|B�ս�ڮ�D�4D��%$�8w����d[v;�;�����i����rpD�~ߧv������-`_�w�F�9��f�"V�� b}F廅���ץAmQs�d��M�~�XfRl��f���^�W�͘g�&T��ck�E��GY���5#B�9�8��OM�̦e܈q��v$s�0Wo��tGϿ��/�~�*�v��������^�y�h�Ug�=���P��Lq��R%C��䏈wp����n�.��S��}��W�q��n�Oq��nǣՊJ:Lm�_壜7lA#,ֱL:�x�|ow�]F�*B3��O���t:��wټ��&��ty!��٥2a�����?3��+���]4e��U�@S���5ƺ*��MR'�w�OArM�%���Ɵ�Rv�?IP�v�7��ꚴصu��B33*Z����v��Cq�H�$�x�٭z���A�}X��k�Z,r��P�E�*�(�S�3 �)����Zxp���%�2h��(�Xy�?F��#�F�N��� ��c��d��g������*�N$>���D����N���x.H�	gkKF�\�s�6�� ����5T1]\�lzױ�Z��Y �����%	,�����."��j�����]ߪ]B"Nr�X������'Hz�?QfD��q��`o��4ۯ�j�V�5ܥ���o6&�ύ/�Z���<(MY�ֳ�>'H��ln*W�-K}�p��PJ�DUOLB�����U���|�r����w�>�W����g�������qIw�P��@Β�Go7~�C6���(iK�2Fk
�{{�\S��.r���2�;D�*F˗*H��=c����"Ձ5qnyG���#W^�GK��|麇Q��Z�Av�V)���SsGu������`��f]�jZ��|�ZM{'�kjI4�5���s%���|�>W*5��bħE��&f�L(39�3��������J�F�D������r]����	�0j��@G`l�A���:]z6�2?4��rc��L:�@�^�I|Q ���Ud�����ljWD��
��gO��n���_Cg��x��?N��M5���%�HL��k�>�N���Ԡ3�
���*�%��q-3%���WPo�~��xq��waR�\����11�&�a'�WG8�6�I� >��P��'�;hP��Vs"5;�=e�r�;L��󄨏ґ|M�V�F��z!&˵Sa�_�+A�Z�YY��g��7I=Ԡ�- �Kk@�0�)_�"�i��]����ѡ���N@i��k;��N�Ģ�5Z}�\8"$n@bR�AB2�5|qiO}QP����u3�ZG�	
B�^1g``Eb�j���F�{�����x�vw>�������ow��VQ0���䞂�Խ;d	y"Ov�r����|JLH9*,gB�?n�7ܫ��Ji��x��&P�cZ�A�<YBOKؖɸ?����- ��O�ϳ|ۼ�w�(?�t��Ȧ��>ֈ|�5��%|�\�x������Ta$���ѓ
���\���Bl��c�3�DȬw�%(A0B:�����(�Vb9��@�,�J��F��r�4f�юI����