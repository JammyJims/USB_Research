XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�@`�l�ė����(�KJ3�O��h[�D�7�a�ŧ��e�� 5���x ΃��ۺDW���,����:�|�hO���>D�|��h������w6[����_�Ҕ8e�)�v[�,���`� �E���%�@�9k:{����O�d�����
 "u���şi�i7��?-n't.%1�y��eYr�I�H�&����fK?+ ���w�c@KAo�`~�qb"B#I��<����KhM6�i/�F�2��[�e�Hk�&#��,�M%�T �PPx��󈐱].�<�1�/dD�5�Q�j��Dk��_�<��։�$Wgɔ�e������ձ�o�e��28b���C(�;�����\�S�:�!��g�����s�q��FU���_��i������.*�������N�:�v]"��	��眉��O��ʊ�;JzKm���+��ڡ6�`���K��_�;�.ȸ%�U[���|����e�,�֬~�ב�I
'��=����a1�åA;���|&XrO����g��Ul}t�����v��價k{i9i��
�u[¨)���t �o��t�k�Kpf�����eյ��A�[��k�u�]��3OL�m)�V�eql�Gة/��2�s��A9k�X��\!��D_V9<p:J��񙘫�8�%���X�NY��C����kD��"�w��g��A�-�r��X&����t|Ӂ9���Ƒ��B�r]uD�?uE��T�'<�_n�ğ���CP�a�_���XlxVHYEB    4241     ec0������/�~׉3K�*��>��S_��ΎM��=�ڕ�3���������H����س<��9&�+�?�z�^�;�#�٬��o4˥�*4��0y��:��ZLr��-�GQ"��;M�UNt���3��~�Ė��H?�/�,�8^�L_⮟\��<d��h��Uا�����w�m����C��hp��x���Y��ZK�o^�٢��^^sDz��# ~3�ٌ�^Es�7�o)#1[F�i�Щ�̂�$���TR���u���
,#1��+�`[�z�E|M8�_ke)Љ�L�c�m�F'����%�hvn��H\TE�d޺��܉s��5L�Z�<����k���5���e?$xu�h�l�._\�4�.����k�y��&Bfe��C�T��m��!�ӷ&e��&4}�X�7�o���Mb@��9�Y9�#���v�^N�\��_U�4�`�B4pk�gX�PM>��c=B�L3��R"PN'���0��}g6�0��+��z[�yȧ�sq
��š���H̅P��%j�E�O3�G��7���I�B�����]�:ĺ&�4G�֌Yq�Te�h�}̜����X�],u.�-6ⵑ5�̆6���~]��\�p�����S�t��?��(����4�w]%h��60�<��	�9n�-�K%��m1O�kq�Ƥ�à_�Xs���ӧ1�k�����<2�Q���ذm25I����+��/=n��a���&%N���#8Q1�O/��Pu��-[�G�� V;�dMN*G���N����c��,�y(rff�<~�Uʝ�ܰ��m����on��	�G�GaEV�s�CP�V�!|7E����-!��;e<|�x��XS��ͦɫ%���+m��L�Rg誘��tk��,OZa���^Э�?>��þ�
G03C���ݯ�s��X�� �"�c�j����!��Qz��/і�%*#"�ŀ.b��YRL
3L�)����&��x�E�M7�_��c�	�WP�$���5�:r����8]�7�o/�)�����񇶭x��n4�sܢ|�O	�"��X���bxm��tcg}9Ƶ| ��(1ڊ��X ��!̷�zi���4��<�l�g��_'��>�I3�Uva�pz�2���9�n[ѯ.�''�-ki�p6J�V���)<�D�M|"O+!� �9�G`).�[!�k�jAnBP��t��fgX�IW��A�g41V �n�G>z��
������Y���f��VB=���
F436�� YA7Ht[�uj\0i];�"#0
ԩ�0� �@�8X:��1�oZ��Jw��H��b��ҟ��_j����U��jWG��Y��;�}^�{n0��m��9zӴ�2�Uq�H�g�@f�TQ�j�*�ڣ �V	?�4r�}$���6(ۃ���LT�yP��V_��E�������[T���3c�*�"$�����7�$��4�Ki%���2�MLZL��iLx�J�D�<hu`���I:��&�C[�=�&K����+�%�jc/V���)A�'��H1����E��z���%z0O�}a���Z:��<�uy��.U!A��J�W����аR�:9�Ѵ$ɓ���RD<�+@�/���5���3ǧ.vh���^HJS}���r9�<��cMS�QN�)��
$:0�n񤱒��	�FRM�ab��;������\�$�X�U�d��K}E]�MP�_?d�|S�	B���I��%���@��޵��S� ��� e �� 
k�Y8I��^8I��˵�C}7^�9^ļ�&}�S�刁����36�_��h�ٜFr:�V�W�,[���؍���s���/g�ԁ���S����I`HI		��x�f����54
���\��8�������
�%����[�o��������L;�w��!�Z@k�#��[9y�Y��Y��`��1�Y�z�^�;�9��E�n��^#F&q*K�<#��LER�2��>���KF,iۭ0 �� ��tCs~EX�<N�GpصVZ�],�lF��1��O�w@� b�Ҥ����T�u�`��Y����?"9�xV�G���n��V}�om/:��>4b�)��(w�sR�#�Х�0C����Y7�z��"i��+�C׹=��'��(֠�1�Dxo;PK�����D�Bvr($5�Z#|�hF�(�v�p�5�jz�~�]ϽzWM�F���J�����{(��`j��D��_Z�>���ꝇ�!�{���+�%!r��8Wj:�4�cPX0<����y0�ڷ��m�8�� ͤj�L���6�hw{�}8�g� �zp����6���RbR�	F;���A�������M��kv}�� ���#�A�XT-�I�I�3�bރ�K�|* "�A��[K
s��=T��3���CJ'p�Ws|ϼ2۟�F��	֖��ϰ!TX��Ӥ�`�:�(��205�I2�ὠ�"�f)>���N���ݴ3��JZ�������E����+~���?2�\X�f��M�G���9O���fVih�OI$TX�[)��t˴�	���;,�dȌ��_�aHV�k�	Z�#>{�#׵ڍV�����D<lE����Ob����\��^�n��ETKS9G���}"�Г�مY�(�=�)?�����]@�c��A��Σ�'�ޙ�B�����_z��m1Ma��A�����Y��q��t$ً��%�����9��$�������+Rx��B�:Z�<�����ݔ��b��Xjy8H?.I;�>�0������ O*��4�� 8^�{��s/:Z�^.d�d�)�9�VEA�5��2�éB���V�/��ݦ�
[���5��8d���0JTZQ��T$
�BL����'L(���'Lz�X�X��gFWJ�X�j[1K���&�ĕX���a?�-*�3��ep���з��$ݿd��l���A����͚��ƍڕ�����Ph�5�Tw��_)�c�+B�t���<�I�ɺ�G �#C}U��b`� ����?�	�����స�8��ģc��?��N�ű�m�i�ϯ؟F9�b��
� *����c���J�N_,��ﳁ���s�/��Vs4���A�Ail@��p��	��Q=-g��R�PV�� �\A�>oy	�A����k�ܟ����:G�e%d��q'��L-!�O�g���r#o��t�{��h,?�E�Y6� ��Ay9|y�7�mp�������K��0��}o����[(�gf�鐼0bC�f�K�Q������'�9�C����1ۭ���^ ��v~�Y�Z��W�J�Q�!J��zHt9�Q�V#R<ˊ�+N	��W�#��PR+G����^����Oh��L�$�a�ǉVg��ߵ��Q���z����ɚp��3k�$�˔ؾ��[iJ�?�;U��H���pX��?�)��ހd�2$����y����K@<�QA�TV{.C(��p'�퀬N�Gif>V->���Y�:��i0l�j&2��o"I�W�Y��rG`d�z��QP����}J�'h��.U�����j��
,ٸмS���6�s�X��٠�����G��J���8�,������S�'*s^r��|_x�z��g�\U}H�w#,�%��{�����(<
ܭ�RL!n40��Z����j}x|�Oi�#T�Dd��&K���`���V�'����9���}'9�V�-ছEZM6�8YO�������R/an�ےs��d�