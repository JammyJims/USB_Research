XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Mө2542`~ej��(�!�EG��������c}T=�H������8�vx�ّ^��m�a��\�SA���#���6��Ļ��L6E�)U7n�[�|-���] ���l����Y�+�U�⻻�����
�~(��ގ��YDd�z(#(�*ĭmU�j��J�#l}~V�y�%�aJO��Zmt\�70�7�QW�ՠ$:}�(�F�a�Q�Y�������Z�Z�E����]�c��2È�5�⇛b��&�Ncd����GSO�������*.�{���	^�wш�-%����f��J�:��4�5���	恚�[ ��	Q����HO�m(���R8z,��H=F˯�%�nØ�P^�Pn���p����bzݾ�/�ރ f���O�K��2b��<��g��K�7,�����2�ɡU�zg�0�7�IŐ�/v��d��x����4�����.܈#zm@R��Yso��̏�� e�X�/�H�&�)m��C��g��Nu�DG�58msE����Ԓk#��0�2Nlj���´����<��'<b�O&ϥ���N�����

��Q[�'���ο�1�ܝ-j\���A<��T�T�o[8�I�����p�IjR�6����-���}���Y1Z\�@*�N�Bi}C�7/=<
l4!��Ol����J�H�`1���7��U.�v���ϼ
�����S��m� ����BdK0�n�<|7w �-<K)������Â�	}� w�5�/�Ɓ�}#�9 ����XlxVHYEB    3855    1000���g�҂TMթh������V���FD>ү��8�.�22n ~.�JX�Ѩ�-�l�[_��� 8m��x��3̒�uT@삑P�[���-^�6��#~ϊ�-�J�y� ���������ii���)�)��@�M<aʔ������c
�ՓW̿~"y����@����.��G�aN?l�e��/������(	�D0n�6f�K���
�?���Wd7@�'S�����˽��bSM�Z?����͙��陗PI�:}�m�ƷԜ��������\
�(�{�9ʗ�9z�ty�=%YF�̍�-���Y=��Β8  Aq�L��ltj��Ѝ�(2�)�����YM�4j�`$��=l�0��ٻ^,�2�-#W��8��EoX
�y�<����*���!���Ƃ�%�v��jk��~|���z��)xΙ0D������L7�.+�X��>|�g���3�)�!��R
ir�h�G��3}���qG�核��s����U�+fH���ë��;(FӴ�zOќ'%[6����wp�w`��)��g��?���`w���kQ�<@�u��2Qs�1;ݥ� 08v��og+ܹс�t�/cD�G�옝g�ѳ��f���
�
a�.��+��6>��X2rS��5��<�P3�x�>�+^����.�"P�Ƥ�b�^0�i��Һl諾���Ӎtf�vU(3�=u��:2�d۹숣�ܛ����W�px:ˇ�V�;�:�M��A�$�[%C�]�^����_�x��[�b�8��;ǜ lG.���9�D[��S��$��<"hN
��� �b��:�𔼮�����>�kqr2���8�k�����?O�
��3̀MiGr���t��V�p+)0�T�`
1��ܷ� �NaJ^�1��ML��DBA+7���J5/K'Q�R]�k�8�R�i����W�ƽ�`e�⊖�! M�$��I�����1���3��ybb!^�q+�՘�<"��y$b]�~L�d�b�R�|b�g����u��&�vYcSY�m��aD��1A�yZO����`HS�Ö*�>�׭W�k���?ڪ�Hh���;I��SVB:��+d�-6�2����*�֫�`I5�X:��B4�1Ly��п�E)3��܊��[^5�|M����F���HxR.Z7,�b�Q�,�fb�T�Q"+��ZOjLj�0�*�l�L5����%��o�΂�NRe=<�N2l�W@Ve`	��ao�n�+�A,/~,�6���$U
�"Vk����ΡxB���|��_c%�*�I7GS��U��:ۄ��1[Xu����[��_� ��H�ӎ,CV�߼z�D5���qO����C��ٮ����M�+�����%�����&>��>/նԙn!�� ��7�����Cu��iqَ�����WL�iԯ�Ԏ�c�	2w�Q��4T��
P�T�d�/�)�(���P
j԰7����o"���^Kмvb �*���� ��;���3*;Cs'��%��Q`�?h#��yP~1�4�冼q�Q��c������R�ɷ�R@{!����a=Ӷ�3o���b\�{r��d�Άd����`�,��Mڟ$�9�̹#�v/�9'�WX''�\���[��� �,MG�˖� �� q�t�q����=��q�z�))��mE�9��ĵ�1�x������z�v�I�m��sኒ��ԉ��s�|AL��f
צ���1�e�O|.AB�n2���l�ь�@��������
��IUN#�A�^�l�t[���T3_����� ���ɛm�<7I�}U��}�uVє/���'�$���)*)�h��?�~�RL45,���oI�e���\jP�_����;�G���dIK2V@�	m�	h���0�12�Պ�x^�s�g�kk!�ßY��`b�o�,^�S��0�3�A�G/s�pNJ���f��Bχ-�
v3���o��+��[���W�$���(k�=ϧsS�iV�3�j�X��1J��tb�נRl��Y�B�=Z��t-;��c�[w=�d\��l͆�2�}p�&����L��_J�8h��z\��������fI�8�������%�E՝��P��(R�X��ka�\X[@�]�X1:ZY���{սN �]�Ӎ%\�̳�g�J��t������IT��/Bm���?�iH8�d��QY��<�V�
x��Ք��O�k����5�p��+5)�4 m��\���<X��䒸7�N����`�+[9�^�ՠƃ�jUnOPE@61b�&�Z�a\'}�i�m�&Ms������'^���7����=y,�E�X�=,,0)GJ��j�H��F
#|vʊf&���^�Q}���E��5�Ɍ� C5�}'mP �L�y���0�T�T�ZE�� U6%�W8�N�Z��2M��燩�d��L�(J�����i3�y7~�vآ�)��?A�-����W\�nh�N~�[�<�9K���FQ�k���ʏ�6�q4Z�M��ֵ.`v��\��ɪh�\ƚ^/
-oR�;�X���p�����@~\,e�މ��	�OF�h��o��;�Ƶ�7�����f� �ύ;N2���]��F
))�n+E&�3�B4|�6���v`o�K���$bf��-�����f-�R�/���ک�*�.t.k�E#�;��dH��IuT��~f�epzx<�Qo[��*3"�w�����s!D�Һ����<�ڈ$`ٟ����N�~�ᖭx�JE|�[���j1�ӈ�5����}�-̶s B��Okϴ�`g>A��/�;<� �Z��]�$���z�j�%�j���4�7& j$;�%p����{sy�~(�l�#o���Y��s�6p������,�|�{cf{��E"�{l~��g꧲�?_���f�FAt���oX���è�Ơ��W���g��9���Q4��G8��R�.�Uw�)�z�K�v.����o�r����k��`����9\�[�D�c��<�k#��)����l�;�b>���
�~~����ʖ��K��z���r,T�. � �I��ٽ���>�x����-�����k0W"�������l'$&\f~����m�sg"��B?�]0�м˲�^��0(\Jѡ�E
"J&�0Tg,�<�����N?��������A����t��5˳��eW�w�('��o|���z�|}�FA�tR��OWo�N?�:�s|f�K���P��,�@��LJH�mP��z��foÝM`����ӻ��TZ=�X]��6��5=�2N�16�Jm�� N�0�*�Q������)&�� �T�%��y�_����*}���ŸҊ>mZ@J�!�������/z���A����%C�N�h���nf�1"n����t��yθ��E�)-��;�%���x�m�0�+�;��2���QK�fί�9���|�O���e Zq� �r*��cW��xϒ� _��@|��J:O�t;�j�j��N�ih�@��{������Z\�NYI�t�J�m�r�n`����}��b�#I�"�/�X���$��J���k#��I�����3�{Ek'G��b/R��b��P\�bՕz���hFe�s���7*-L0�րD���Q"M���M���
�/�Z:{Y���ယ�\���mB�T��`���f�Z@�RN�eX��CQ�=���n@F��,��qN�t�9�H� ʧ�����?g:�B�6�nʈ�!b�d��+
�'�f�&(����)�r�k�m�b!NM���G�]��ԅ�^[e%�Zҷ]�����g
M_���}�k�	'��^���q��2�֮N�S<������$L}I����n�r�O6Q���#Ϣ�f�U��,{�k�/�|9#c,�[2�e�Gի�� �
J4'!l.��`���>/�͑%M ]A��8���[��2΃�j�Bp�_d�6�ʾ�
W~�h��|:����ܱ�ۆ�I� [�jQ�O��E���;�ҨQ���(�+� 
0����~�%
�ʊӁ�E|����W����9�Q�>:�O�n)����/I�OiP9���Ɖj�v�_DG��Z����,�*b�bqHǔB�vE� 