XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���sv��8�K�V��7��!��ѳ���v뛯��%i��LC�{`�E�{8�ɠ�V�dz	�a����@���O��`��W���Ɋ�β��T��q&H��������N��w�H���M�qRL�xX�F�+f`�xC��6��$&��%��U����^��˟	c��3�U'X�Ih� )}�=ꍭcNݩ�(�!2�XQ6p��@=+H��0��!O�J���3�>�mFT��yu�޼ypp8����|Tq�p	��ݥO�Anv�q��ˑ��YAZ���z?}�fl�7f�`�ٜ��]J�	�!N�R��n㇩�V޵��+��|��>���-#��p� K�L�����ȟ��;R.��1�ɁR�-�$�+��s��y��K�A]����$+Iꅯý�ۏ�~DM��5n��*d���8>����N����A�)���/hq;����D�kM��H=D�B�������B��7�.�Z'��H���k>8q�����+Mo�<�쑗����<sB���Q��T�����L�
Ҕ�0>B�S,d�cuuy}�[�Z� ��l�d���c@|K�lϨQ��X,�_�,��$��L;$+D��"�f����pp�����A$c�j	�'
�fڍ�B�-�z00�X� JI]`�6z\��c���|��{�!T�zƹF፩����� ���fUp��VE���@xR^ş�Vˀ�<!�̀Q� ��i��$�`
~LI!�FW�4Q�~�.Wx��)H%�+XlxVHYEB    3db5     d80.���H޿*��]��قc'������|A�gˤd���~�nҸ���Uf+��dA4�}�AS=$ҟD:�ua&�h�>;v���FA�/��C�M,� v�_8�=od��S;�_�6���S�;3��q��q�M��o�����^����3���ð���~��΍(ï�&�e(*T~%�]�~����p.��,��(o���,�a.-~\���z�XYR������ݺ>�Nb�}K�V�*����v�K�ǯ'%'ux�;idB����!bU�6��h����@Dm��f���a��i����}6q�S���do'��� Qq�4y�#"Uc��|����t��Q<��ʢ�ݯ/{ٔ�>�=Bcb֨�� SϭPh��R�-Ǔ5=/�����43^s�q��s��ԏ�*l3b�SM>L�]o��M�l��S
���	����nG��Gڦ.h��t�O,ND
��U�A
RK �`�$LҬ�I�T�"(�����ф��H��J���LGh�?w�=X��Cp������5,���q���(D�����wħ�x��?
ڔc��)���Jqvmd��Hj�����7r܌�]th#�o���k�Y���GY^V5R!�=j��)/\�;�lHNJ����D��W4�;i�^&J٭/&��;Uw/�o�Xvs�%�qⴂn�TD�1��Z����.+�[��iZ�4�xpq�Ne���#h-����W���7��6�4��4�W��V>Q|@Dh���Q��i���B�)ˌ*$6ڵ�ăT��WH�Y:cu����&|_�?�!�Ŷxh(���f���+"��B���`�P� ��k ��ѽ�R�r�+\3�ʫl���W296w���l!���7�%vM����x�¦�YoĂ�Fݚ6Gbn]bz���0R_U�UK�֖#5��$ɦr���4��0��NdJ ���J��Y�t�u�'�ْڃy�e7>@	|	ct3�����M'^0�A���9�7��
ڶ8�����v��ӊ�>��
�P��{���๕�ز0�Bn%��N�J8���o&,W�j�hS�InA�T��(��G�{t�G��w��>�W�m7����xf�} ���zoϞ 4�$�$:`̳wF����)�����)�P��e�Ϭ�t����bw�mD���8Ӏh�EU8�O�7����#믞���F��Q`P�����.mU���Hڶ3�n�AW&�����lRr����B�O9����x��,�Y�-o��(���?3�7Ƙa� �������Ȼm���UI������J:B"����U.W�"�ɵf~	4i�n�!�X�jvȲ�����7=-�s��%��T	ҁIi�=ðћ�A�����'(�MB�#F�!{�
����jo�QNr��u���	3ʨ��E���L�`��poؑr[�^8Q�w�J5YH����>hr��ӈ�&��?e��$ѯ��V�)�x��پ٭hR���0�t�!��*��m�b,9��d'�r���? �zl�@�9�P�y&��~�O��a��-1�$��<D��hY4x�h�.�a�C�+�S��TQb�BƗj*��U7��c�8ں����+�\yGl�R�ܡ/�Z|ĩ���re�.�L�sV]~P]R���po�t��|�""��j-�[����� �\_t_4&��#R�5k���y'{ 禺H��7�r�N~�y��<�u�$��O)��YՋŎ5�6)��u�֭(G^��#NYޣ��#z+�85��>f�3^�V��p������x��@=kZO� ?^-
�e�ǅ.���_�(��k܁��vH �^�SJ@��0Э�-�䅚����]Q�p��S��g�D�� u�c�XN=�g�d\�$����?��!�ȡ�N@��UŃ'+eby�0�ʯ��7 C(Ndc}[��$(Ғۄ.N�T��=a4��׷N�������|v;�W!�=# B�'����k�j��I���G����s��@����wTW� �/���F�j�=��k��.�q7D��#��[^֞o���w-p��$G�@M׺@u��}��	L�P�7�<�f�^Әs���0M�egaՉ�ؒ��Q>�v	��:�K���(�	~1� �'�v~^wS�v� \*�%���bEx aִ��J	�<0l�3���O_�R}�.w����I�!�d�Z#wn&1���{��K$ 1~i�'x�H�,�߄�/U��w�N��<9�1��,�գ���9ZV��bݢ��.gN��k��iN�DN��@S�Olc"u�'��6W��9D�P�6폜����7�So<��f�G�'��QX/mw(��뻅ޟ���0zՅy��L��A�m�E<���®�ݱ������K�9���ʩ��=��=�Lu�1_�"{L��k՘� �4#�6�N��΢�ʝiT?俲�g ��`����,�����Б��2��I�J�6�R���L��9�]6�/�˕�i;�A�@�t��S�a�M_������Qv��3ۯ�g3���LGDp�>J;3�o�^�ƔGv�*YLJs�A�5'��W�c�3�9�_ul�J���e�^�'�̍�K	� ��&T��/��&�!�ȣ�{�����W4~sJ��g����\U��\�1e|DFR�`��,h�E>�*cq���� ��$lTD�`�6M�,6(�2�n�ZKN�"�*d��v�#0m��$^͠����{���T]�4D��F5a�FB��\6�U��W�am��6��W��&5�ЪB�4�����5�I��n�B�t5�P����-E��"� r7c�u��2SwFb�i����`Za�أ�Q�%�A������ikq�+�v�r���|rsO6�۵��z��;Z�u�3��D��Xv�+y����Dԗp���3�82̐t��*ް�R"	�E��!e��³.>��q���������vv�5��ٙg�*w����M���QH����&S�
U3''����WR&%�,u�G%4 i*:Y������.à�	ڽ��zy�W���_]�v[�lA�s&� �V�go{�b�����0��9�Yt��heU��y?��Pd-{I$WTj�P\4�������7�яxr{�Y�W+F��{��5���� ��7���8�L�c����8����@Ư�%��GK�͡�n�.���$�ƝU�(DT�(�6ߚr���>i�b�vF������>�ԈX%v�ܲҌW�"�Ԏ��K���	�_,D~�\QJ7�<<�8�Ռ�r~8%=�-��e��KE��M�Ss��~na�L�ֆE�	 H��s��T��:́�ǳ�X8Ț`����������6�y�5�)f�M�Q̸"#�K��m�4�J�M~��e�9c�+�D^