XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[G��;ަ!�|�J�e���u�����	�_"o9�p�ms��vZ�F%Y�����2A�b��N 0��e�� z/�r�Gr��HI O=��N�
b`�k�����Ղ>��X�rf����h'F�,|?En�B��jo!�4>�{4�,�П�����K*�+Bi��H��.��x�Sg(�"l���s�K���׼�.�FY�ݗ1�W�g}���£A�2>� IH�� ���VЈU��)�F�R�BrKn�*	6�Ox�l�D�nQz �<�~���M���,����u �":jG�8�Q�.�]�0�����X�b��ô�#��w+��	� �����\�{B������Q��ít&ܱE� Yf#k>1)��=�n��]
�bd��=|C75�p��gcR�J�G�|�2��'�f@>V��i�D'2�Z]�t����dւ�^�{��K��|LȠ��ȅxi =d���U�g�eƓv�dyh��L��6��*�^`)��]`�\�Cd��}Oy������S]�X��N�Eq�Oո��Y#�W�$E�f�O��x�M�}g��B��;+;�r3�@�a����^�>tD��#.�����{T���F������ݗ�X��� A����f"�=#>[�U�5IAd����T��ڏ:fX��@��<�=�"�`mW�֠}�'�=@T�ˢH�b��Zv��G�1���w~�� O2r�[����4�
+����m��ZaBu4M'p#��XlxVHYEB    1552     790���!��d��o���b'� �,����v�]x�p�s�w��{�_����N��k���)]�	���{O��	��
M�Z�߱�Yܧ���^���
��p>���;�!����9����xk��*�+�դC����V�rҲ�1�!�j%�,v?���v0aj�Q�ոU��?�*}���Ů������n�x����=ŗZ;Q8�ӓ��\�|k���.�Xr׎��o�2	C�'"�j�.��0qk����S�'�M�����ػe$�� �<��2�����GI�96�ͥ��)���-��N`g#�TdB%�T�������h�z�/��`e7k��y���{��м� J��|^ݞfKҖ�D��λ���W�`�7�Zn)^c�{#$4fA�r�Z4W�'���Nz
*���v�,��z�l	�	��h�f;����Tԩ��魥�χ�si7ġH�1)����"��ɘ��]�r�[�/6b{F�z��E�t�$�L��>d����+�?qD ��/|�{k���ET��S�sJ��nvRU��'�gT!#|b�{��H�*��K�~��l��W/o\T��'0�[X���P~���8>&�i�R��)�C�����U�4֎�dA�m��Le�K&�Dm��_��D?�8�p�*)j4�M	3�!�ڃZ)N�Җˮ?S����:/��i�	�P����ST�	�	��?x�r�7���0���
�9�$��F�ό�d������f��2����_�T-կ��Wa>����x=n�(�7X�@�����R���i��Zw�񹇥�Qa��e��P�%e�WQVsm�������ǔ8���^!����ߩ������m��v�yM�{dED�	h��HծL��1w��$���Uv���aC��%R��J'��h�Պ���<�&9=��ڷw3�b�0J%��y��� ��M�/9��������e�{���>֊��w�O	?]87_KG>�B�[sK ꓴ�0�Μ�hH<h���돽�����"7Jk�X�|I����9���=���q�"���/E�]�Bza<��e�IH'�v\��^h���ea6Z�ص�� �E�����n3��hn�&�C�\��R��W����6U4�9�c�S�l�"��"��R��7��U4{j\q��=T�O��X�"��Pr��AD�J��̡vI�����z
s"��Ԣ��J�b��}5��ǿ௤ÈK��3.�0df�#���9��y�_����#+�tH�H��7�˹�ٳ�cũÌ?��1�����6~��v��ɞ>v ey�<3�O��I�ƨf��Fv���n�~
�����!���Ԭ�1m(����g���Ѝ��ʶI�W[��A�7S����PX�6��Ɲ/���e����GW�	D�b:T���h
���l����Jx�{�(�e�|&�U��nq@ 9��#ǆ�]�2R�S�^�.�H)����Vy����Q���~�FQ�/�������?YHÐ�Wez��j4m�8��*ūV���+�}�4%J��_� f����ݖu�5.Qݤ�qI���OL�8�3�/[*���XBq���V�g������(�R���wgh��v�[�ArcV[��l���=41�mv/����'��GP��#w��(s����#r�3Pu�j9��$,���t�6�I���h��z�����_ogiS���ʌx�Y��P@����*t,�o����A����0ھ9�Ȱ׺��Ƈ����y�A��I{��H���]/��ُ܌qӉZ���S���&1��@��< 5IN�&�����|QP��G0;�r�}���gN��T<d�/��P��ݚ2�M%DF 柰ѬN���9���X��0G�������n���Ww��"��c7* �ot�ɵZ�]�[�-ﮍ�d)#�