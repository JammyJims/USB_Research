XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͘��}���)v�����lU����J�k��`C�������x6aq�Ʃ�:[u*�V��=>�����=$�f*�wL\��wz�6 R�O5�ݙݙ�"Zi��?�<��)�7�:�6�g'~������n(�[�c�kC�j�Y�u�0=��ˊ��A'�Aki'�r���l�PetWz*���V[Z��c�����c:���L���Е�'&�i޷��KvV*jo�T�p�"-�y+��@t�V�����ZL��5��|	ϙ�5=^��Mq�KH���a���4����ݜ=fz�v�Y��m�?1�N�A`���"J�L��[\_E�`�#óAo�z ���8U�X}N4�����}�{ːąJPܣE����R�3#� ��E��wP�Ѡc,���8�>
�A1 uB;N�������2^q����s�#�$�M$V��UPƒ�K��I�d��[�8[ �!&�X0}q#�K>��"R�`6������p�uonh���s�`E-{땼vnԺ	X�#���8Ā;�W�V�E����+E¤p��ͫF�¢������~�)j8�F�H�8���x	�	&F,��R4�~ywhm������.m\��T~2#W-�U�>&�]�)o��>?�R����T��U����5��T"ɷqR����RY��9��xs|�+�&�X'�!_;����v�;\���*�4p�md�Jdj�8�����`���c�CH�/��?ȷl킜��O�6��nP'�7bi`۴�	]�ZVXlxVHYEB    fa00    21c0okE3��Xj�*:k)p���ٜ0v��>�-E��\^>04���M�$^���p�_}*���������Z(^����!����)�*�6��\��`���Il���s��~%f�|ZJ������(��7�pw~� ��n쉫�̿!���N��Lz6���� ��q�$�����4�k�VU�L�Sۀ��;a �Β��6o$m8�}�5vE<Ȫ��2[�j�z��j��V<!�؅~�k�z�`�j_o4�Tu�����<r#�8Z�-��8|1�d��	q]�P���3�f4̡e�>fJ�i����������Z��B-�d-��ʒՍC(A��?�����N�g�38����
L�7�Drw~��y&��˂�	�Z��N�U4�
<+�Ԏ*�:�y�C�j<!U,8�\j	l�_��+���4��hpf.����_ �&@�W�\��:E2��a��G�8y)��w81	��9�Ui�.�>�j�Qe��P�0��ɼ���g~۳,�f�l#��ǻ�tj��ٙ9C����q0m�c�E�n���;����,�� �o��b>�vb�+��!I�P�]�f��ߜS�}�3��n��Cj�� �'7sc��k3,�+6GS�-��fq�͸1�7��B0>(��7`Md�=#�'i�M��'��`V��X%w*j����06(恵��Z<��(Y�ۻg2�f�Y;�yF'T�X���kF�X��6�H���	�{Q�T�)�	PJ�LF�ǘ	tΘe��,��y?�8�����@u�lc���?���sڑz$%�Wbv,�t���D��:�\�W�oF��~<��c�.�v?���"��Q[|�Dx+�h��Xa�v�M��2�35��s����L�;��y��L��(vb;q˫�w�K�?dv2�T�[�#�W�0�]G����d6o��!2Dy&ud�_Am���\#ӎ��X�I���pEo<{UEs�X]�e��[�'L��:�:�����<�3x j��u�w�<R�_И�+���=��9��d�:���[�i��<6��eT��A�H	� ����TEd�{Y�5C���qɩs�*@��$:ys���gF����yNA��+��|��{T�׉��=�����LQ��ǩKh������r
��	w���:����3�Z=�wU:���o,�b~�iױF�k�����Z$cvN��w�x�dg4,�ƞCs����\�5m:�s��i2'��3�ꆐ�s�Kvf1����G�c:�m8����(A�	�r>�`D��Dx7N�-Z�|�<D_y▦8��{qG��}�j���"� ��*��(��b��5��pz�*��eX��hLfL���w��u�!��n�Fm�g�;%�*�&lU�F�v+%iz�&���;!]v�\"'��O��2Vp�3�ܤ�+Ŀ+�t l�e��u;����,8y/uJ��~�,�Um-�3�"���w�`$����*�@,�+��{�f׊�G�#?ɯ4����a�X����r�M	1RK��I��+%�H�X����n<N�ɠ3{-�����2y4�B�6�2̩AN��H��!�ܭ�5% пe����vR6�ɺw����f.�N���A"��ո�t:ݤ�{Q�+��V�7A�l��� ɘ�[.�'�wNN��&���V��m� ��5c�@��|�}t��U��!�E�x5r�8��e�P������[��׆��R5�߳��\���ԛ^Xq�㿙W/R������Q��{���΢W0Hv����#�P >|�ڮ�_��<��g�b�u���j,Y�AM+�9b1vp|��We�=sk�s$Z/�XE�Ӱ��et����o�('CW�� �N�5 ���Z�^�L�h+̗�cjU���[���ZA!$I�6ߓ a!)Y$w{h�U?g`o9�g g�:������d�����4���|^��q@؝F��R�)ʖ�k^p�P*r��A��WA7���O��DC��)��grN�rś�	�l���D���8��m�j@;�:���{m�&�L2A77��!v���i��ѰO��h]�Y�,!�T�:�īO����Ui8"�5_T�:4f@6���I2Pݚe���	[&U���Ṅծ��� 4�s����`1�J�8|r��S���j?���+&��_�7>2o�פ^��j ���Y^�_�cu�}�̶�s0&^Z������I(�`P��AL�5ݏc��g�����zh�H��ZtO%�;����^�-Y�S\�Kw���l[)�t.3�'x�
<�!d��i����<����!��|���.2O��ntL�Z��x[�C��N]P%/�Y�a$�nQA�'Ed_�%oUւ-��{�
�4������O"{L�v�/��7K��.�<���/��d��#�!8�M������vƨz��'��Ք�`G�g��X��[6Hw�&2��gΥY#E�A��B<3xE��U�,�Ì�үqL�o�����w�я������W4�P���� )1{�/5�Q��"P����8Z�x>��[nk�r�C��
	T���<1U��ڊ�`\��L��0�UR�Q�(R���>���hPN��_6��$Z�ѵ�ȅ��^��aE��� ��4��ّ\�ע���RT���d?�T!�1��e\t~�s-�_��o��5���4�'^Ly��S��Ka,#���p���e��B���k��5��ù+9@"���~��K`�a$�X��n�m=_����f�
�k�ޜ�wBHH/VZ�c��M��~�gV�w��b!1�QL4�`����f�N�� �GK���eKϞ��@r4�q�c֥��((E����
ێ�j�M_��b"�����肤�f�b�m��(�ݙ�>�ԂM�g�8�L�(�i���+�#���;��&	%�sBa�]�5�_dq,'�,��v�u�N�8�|SP��hc���ݹ3T<X����>>��=<�����M��O�R�G�Xj�C����*�**N*�+:{M���S���ϧ��K���&<"q��u���¡覒�����d�9�G�y��	�l��h䐺�����5�&'PS�N��
������/E�z8������8����:��enX�S�x�*:g�����~��8v�����T�:�Y��A�g���w��	�r�wz�`���9v.�������{\10�=u� ��֍BS˴����]%#n�������Z���*����0�����PW��o:���~�e㜥@���~Ȩ-z����oX{�_$��1�2�.£:ٕ�Ms�W��vB�kW��#���+�����Ԉ�p����P�w?摒�������(R#����F���iIc�g��dSŔ������
���~0ȁA\�/�4jZ*"��9�0������g[���ƹ1֙�ş�5u��iA���5��h	=-k��W��`j����=�"�"��T+����GL����~�.��-��2:�/��<K����rף��D�[�A/��2��`�߱�������������(�~���4�s�E���m���8�Y2|Pcl��3D�\*@�H�c�&C��Mk� t����������jटA6Am >�~�/g�Ѿ�/mD�U��ҷ���m*�xJ���QGV�G��'��v��4)5~&�`��H�[����+�zJ�P�YeZ ��Õv�C���@>h)40"�&��ȥb�@�V�o�';��58� ]?5��U=�)PW��h�� �&��^�d��+����:��e��uf1���A�mg|��n\M
9So�wu;��"�*l�b��+�[���G�����[���F�y���/b�0�q�����;�;wX��*��B��6���7�YH�>T�)h�s]�\x�
�0�eĉ�pe�pQd������{t��A"�o��W�OG:�ӌ��c�7@ZAx�����Ę����˗�a�V��p�Rr��2|ꬖ�z�ӄx��0�|�ڈ��4�ǵ�xfd�#|��\ �G0u_t(!�����5t)҈)��Nѩ�4]�
���J������_�z�L�Cd.W�����L��m�U��j��Y�;�Fn�R<9W��p~��@Y��d�4O�ߨ�h�i��b�5��DZ��ү�趏��r�%~5�^�"M������oJ×�=��5(Q_d����mif�-@���x�P�U��v�TU��{!=,�����x�^T�q{�֕4[�R�uoT�0���I��1�0���^��7C8���G��B�8�Fsΰ���lfa�B6o����#�j2�%M0�GKm���|��tPeǕ�Զ���㌸���Ν��p�	��:
�$�R��ձ2�&d*.09Ac��d���)���7��4�xY��-�ԋ��B"�2�\�K��F�r�=f���|ERP(��*<�T��@K�������1UwT��sUFR�Z�_y7�D\���*R���2~��TN��j�jN��*���w"alIt2�����yw��\S�;�9��J�m�
3��'�Z�'yK�0ښ��ކc!�kLZJ ψ>@@)ް���
����<��yaӎS~�y&
����	�[Y��w��h�%����r����x��� �c.|`�aD�H�ys%��Fž��XP��(
������=l�3���Or�]�j��F�2�������Di��?���o<W�e�>F��C��c�"�E�IS�x���{O�ᗽ���u�\(JȴK���/�:�$��k� 7��A%�Bړ,>���$��J���j���(���A6� c/w� ������3l���5s*�ks����=B�������0`_t��?���+0F� *:� ��;j����_�{<3��*�a��~�\Z��'7Akl`%3��������c鹨��CR���o�}<�g/�g���3����"�ða� ��Q���CwZ�Bz��Eg60�JYɬ�^?����^�SJʷ�#��y�Yu`j��A�;#uk��������Օ��A��U���3�G��#���J����lv���|"�T}xl����%;�Y'\�<�4�� ����?S=�0��x�s	��{�>��<�x��t\�߯���up;�0�~�%������R&�����YpH�1��DR�����w�G%�Q�1b3���viP��2�o/~o�(�v,s��s_�*F�K��R�2�H.k��B��9mv���ͅ,N��pN�y������=�ؼz�ޗ?��5�ڲ��a�1�d<=�~j���A��'���>�1�{�i�m?������^��*y��h4�^��tvINZb���c�n�xa�7`͘i��	��PS�PFZ<��sdNtY#�k)�_U��6b��͌��a9��G˰�43>��D��O<�P�>�=�c��b����k���$FG�D��
.�s�G�����;ٲ5R �|Ȱ�&���_�e�m���c>ճ{�t=?�zC�I�09� �<ਸrMsj��pF��#l��GŪ�Y>t�W#��g�N"�^�Eb9���yE�"tSx�eU�c�_�Ӕu�.����je��-ɛ�$�����C���s��=��TQ��&�8��Ž��:�X?k)�U�lW��N�1p7ҡ�E1O7t��٢�U�q�/{���Ⱥ����O\ q,����
9]+��d� ��*�~wb���G_��KB�E"��:R��Q������ı�1j&�Zr�.V�.� �2O;����1�n
3�Y#�Y.`�׃�����s�)�Yi.C����ӽ�=�o��(��O�0��H�}=˙���ԝ$��`c3k��[�V}���� !�{�#���K~�K�~���	j:��s��כ�-��;�P�̶��C�>�tw�*�rU@u��a���b�~ލ����ٚ<;�H�OE�ꍲ݆�ҴǬ��u)+a�9���S�^�޵���c&�,>#,�����أ|�uN�w2Z��CA�o,�~��{-��������Z�d�@�V:��� G��6�̺�W�K��>_@#=�=�LH����߶Wf���z.�ϖ�yLW-�������8��i�U�b�� ăd�A�"V�"�n�!���h�GŶ�;�aM��{S����w89���wD����`�H��M��-p�2U�;�\�x&r��Mb�A��X��hn�|�*��>����O��'V�U>K�Y.��A��[?H�7"����K��\jͷ;�~�4�Og�@Fn�7��Jc��F����4N�z�WT����������|��u"|��Q�N�6��R!N'X]�'D����"��K�r����Z�\+�t�8��bJ����=uZ����>JemÍJ����B%�����I��~�u�זͷ��e]1��)�H:(�3Z��"��	�`����ڈuhe�m�ueyH@��r�����܏�G� �����j+T
o�ؓzN46)��)�N>Q�=-Vs�
yh t"���ǋN���_(�愵~�2ԝ�'���-Y3�N}B�<{�
��'��%�pKg-0=��JQ#ox��ca�&p�ܽV�{�n�8���I��@�U���无�c�\�� e�Zr6[��><�fV���	�6���F�p- �yKwfV�}3�
T��䨰l����J����M<���	b1�-ҙ{�)�ͻQ�T7V��q�v����>�	��W|�b/!�[cRB�ǿ̕o��h[�W�'�����kcU���Y�w-<�ߐa�ު���`ݢ����n�;�*�\z~�ģ�
ܵ�e�1�H�JuE�����Sui~�4�T��b����lu�D� 5Ȏ��m��al%�O��G���:�� ����Kw�ۼ��o��H�dB v��xYp��"���)
�|g�;Q���E�X���~Ч����]�]��������~����z�����;p�3��Di ����A�y��
=��0���$��.��@��"9Q��wV���o�RNgsu"=����D���ҠJ�q�Ӟ��<���lT��"���:R6��{n��k�{�LK���~s'��\�M}C�2�/�">(��j�Z�.���;����F�E= �M#��TL��5�&9����;��0��y�9�UZ�'4_��m��6]t��k)��M
�e1�F���o�b�cnl����a*q�文�!����4�_�,�x����������;�pѤ���{�����F��~��~���L���5e.�Oޭ�#&�K��N��I�_~�5Qi��Fj!�ex=i��̈!�hE����[+��Kt�u��(>�g�y�6�6�^�NfK��y���]��N�ep���[f}����m��5�2���ưw'��HGo���y�M��{��1WH�=.�X5�ɢ6�H'٬��>��{L�w�0N�,^�X�5S8uߞi>Ο�Q��<�����o�Uk�fJ�O���N�����Y������G_��F�;�L��+4��^�#��|>�a|0Q�~.��5�Am�ⓚ�3��FVI�=���]PCn�s\0cT(R�=J�[��k	ks;�M`�eĭ&��{;,���Jbi�c8ӄ6��*+�n�%��UmcG!�9f�f�B 1����6҇c;Y��� �.2�wdr7�Z8M����[�r{���8�p��$���1)��`�~�c����f�bu�� �.���Y'Zn���� v�TpC
�T�=|Yw�;H���ߗ>ѼJ�=�E�?�|t�n��Is3]��L�Q}X���_���ɞz<t&d6C�<%�{r���~����'���!�S��[<P-�UY���Ǐ=��Hl?�R�_"(I�ή��]L�@d]�C���.����)	��o/���4lŠG�r0��&2-3�!�:yR��I�%d��Ux��ئ�1�ކ���(�۾߽�_�zx}��VMR��H�S�������gWi�Wܭ��L_��gѦ%GX
����H^����DU�N)�-��%y����IE�(�����3��ٱ]AT[5��0;�� �|��2��z��>'�6��zP�(�lN�D����8�'���$V}�I�XP�;�:�\�[���2���±����#JM��j޶kߛ��cy�z?��z�Lҋ��`��R�w�'+������٪<9�l�@�݉�ŹI�}t��幭���h�����t�\!#�DIg�!(V0�Ҵ�XHm�:�ZL8��2��q�JC󽻅Lh9��:�|����k��a��*�t��ۨ�)ڥ�SЅ��Á����Ҹ��\[{�=T��ԯ#�"�_��)1𧣚��Ք[Zi��j-Z'��9j�����nZ,��)��e�[��l�."��~0G�F~��u���՛G\���Zo�{
|\�0������ueFί'<�pz�)r���;��� ��[��H%I�pg���<D���·�T�s���G��t�z���� ;�Iّ���h�:8Q��lF�9ǣ-㻛��@��ɑ�cX��Hk���,�?�m��ŗ)H#�f
�	Yz�؜XlxVHYEB    2997     720B����.
��|�3���T�,?��>�?�!AG�ְ�rC�&�'u� @�?Q#-���+�pE�`�hE/�ZV*	�����7��L��Ě@ަ�'�j��^w�y�����n�������,tⰣ �3�E(pȬ,��A�TK&�|�ٍ�{�Ų�ߵ�X3�2�%(^�^�K��K|� ����"�OX�7"b�ڳ&�F-iޣ�`p�C��fe7���]�o]�N�j�%ޠ��^]W��j�Z�Q6�9E�Z���[Ц<.�R��!��ƀ���:g��V"ȥ���"U��+^��7�"��¥ ��'�C� �`��K�Z<ҪE�&T���xyw��(��޽x��#���^�h�/qqx�ʵ�"]8�6��W��ֵ?~��Wc2~��N6[����7��G��a#�3�_�X7J��j�E�J��5pF�� �3�9?�6?R	��ew�|Jlvѫ��s�Pۚ���/����m�C�M��=���1lw�B�[ |#�?(N�5��/c��
����p>���e���-���Y���:MR�<���9>p����Tw�۞���RKm�ٕ�W}�s��+���n�X�v��q�n `c�Q�⿎~��LT�^xPi	:Už����P�t�����B.ɩc��;�,nQ�Y��k����"ԈMtȝז��(�lAK��HC�x�Ep�1��ݦgA�y6=��6��	H|y9Pq�x�����.Da�>?#��M�����ߍ�NGHi��LC!"0G�\��q�/�^�.r�[���Q.�e����o�Z�<���ZӬMF*1g���i����E�������|R1Ʒ�
fC�C��?�>F�w��w�y�9>�8~��$�h�������c'G�{�y�;O�`�����J�o��HZ���8פܐ�Y���J�'.o޽AA������]O5J����(������e�������>�i������Y�W��?�M����^4	���p����4������[깹W�&�� ��pt~9U��T��i����v�^Gb�9�][��?�|��W}��+:21~5�4O	]��#:6F�������ثNz��7`�q�D�:`΋_�sx��fg-���-@�tW.`�HY�Yi��Ղ������N�q�RRä��37��Eud�$}��`��:�v�8d��1ƍ��ա���E��5W�[��̕��u�W�z���³<��G���;
P �0�/���#WJ�=��P@P&�T��\[`�%��3�5x ��ӥMக�*)n�[��};�������aM�yj���ƻ��:NWA��4�;�0�b�1Z�br��mskQcBdW�$���~��&U0W�F#��Ӻ�^SW��[�u��@�8� >�7�~�K.��IR{��%��^|)�AfW~BY�+�ھ����N� ���T@
>�����o��Q�!�!�g=<$*Zf cE@=���l_��-�ހ�G��[eh(�����>"d���Tϵ�'�֜1�o�zx���}�_1-e.e\@��ɋq�+�A�U�l4z���~ơ�)P���$����X7�� ����B�Ŗ0X�jȤ�1��[�rGjtk���y�%/�1��k*���-H��y�Z��R@�Jx4�^�a�����ͺ�]Nt'�;�!S@EQ��K�a����H��),AX�0��Б���	�}1v�T�Q]����ǂӦ�x��X�7+&�bܟD2H������]�1�Ea��pfP�e���z�X����qi��@T���&v�rp��F��6�֚��mH,q(�����q!nٗ