XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m��;�&�(��`֓�d��+7ο�قk@��62�1��K�P��������Ak�D��X�f�3�gè:F��cP����2�GXw�ݓa)��DԻ��p�����j�a 1���	�|��hY�F�r6��$S��u�Eی����f�-l�)΁�c�h2F��r��p��Y-a���_���U��-�:(=EBt����!�7�W 1Z���rea�G:]6@ƾ����~�"�؃*}�`��T(�����������t�?���Xe����ػ��pj:�H�=���昀�h�-��	���Kr6�wk�����qC�05dW��j~G'&�5�RB�(�6�D���"����ql��z��������ͱ�P��!�P�8	��H���k�x֗&�~F��az�2�-��פ��e9w[ �e
���0���x�6����p�8N���z:�J�&��°MK|���pYD�CJF�$���p�C�_�U���8y4x��
�*�X�D�J�Ǖ��}S����Р��@��ǚׯ#R�g���Y�W���Zg��h�>�9P�KuW )�W~E
ZѤ��:���R�)�dyg�z�8�s�h���Q�{����`�&��$6Kn���" 6'��\JW�|��64z[2L"np��Y���1�\�'���B��f�°ݸ@�s�P1Op3����sο]',�����t0�f�:���ꞕAs�м3Ӊ�E��ן|p�Y�l���~�	�D���Z&�?�#XlxVHYEB    2bfa     e20^i��F�;i��ν�ʛ��w�]Ai��Vv�Τ�a.+-$S����{H�㒬Fz)�E!��4�����(�H�jA��5�t����W`W*6ٲ%�I�ͤ����yf;r�M���j	���\�I����^��b��,&�w�aS3��m����J�:�n���T@%�6��S(�Q��e,}��dN���?��wԘ�Ԛ��S����Q,ŉpRWQ~�kQ�AkJ��-��l
����ψV˱�VL��N#i|	���ў����[���qb���x8��+tc����J�ٙ-��+��s��/{Mԯ�����t��Z�����+]+���[�d��H}��i!W��M{�|e�Y-�
�� ��,Ҡ�j��ͯ�1������#;�]��P	��?������>�ϐW	W�$,ϔ${�qd�"�KZ0�]�5e�;��(][�,���e6�vb�5�~���� �Tu��	��$�B3�#]����z��#/�-p=w��Rd�;�K8�������2���}0*����CP>#�;����rUߔY.������3�y���~��6̮D��sх�b����{%���6�0\��	�+����%�O���A�Z�n~`�RL����D�������@~�f��Bb�s��2�3]��������	�x��L-s�t�� ���7����+�:'�j'O1���>�A��;�S�V{���=ۂAR��H�����0�c`�ą�D�{&��/d�ХSX���8���Vtg4�����p���~<xچ�Ɂ��l�Y���|��|=+e�>�qg@�C�b�I޳���r��m�7�m#�Kxl�/��ޫWЊ.|
�6
���>����bC0J�d{����m�rObkE*w��{K��?�߮�=�r+��b@��$�a$��,���LŨ0��>M9J�ы��	" �8�q~��|�aԲ��#C���i*�+�=�D����P)��W&.��Z���a��MK�������g������(��q�	d�Y=���$_z���'A�+D��C�gѿ��T�K�z�>#�#g��Œh��yǪ��J�@%�:�^�No�r������ux�cG��<En���]/4:6\��s��;Ir�}"����]W��A��Gy��ayyZ
^Db[�g:�I&.
�!����HAu�ܶ�d"��ݕU�C��h��M^xa�3�,L�͎ߧԌ�<���rʸ�yF����AR<tT�K8s����xd"�Ҝ {+��/ȴڗ/��҃BF�/k�������õ=�_�F�OQ�L���-f\��"	�M۵k�О��-��#i 056t�y��0��O���[ɲ	�m����F	�����
烺�b���	!�E����]�Z4�d�[�)��M��tg�h�x^R��ј-��� �S�a��EK5i0��� ؠ��i��S����6�~������5 qO��v���SX��3�M]�4���*���E��͈���S�i�s���/��p�8�)`Y��Г8�-�:���WpC��7�VR�&9���9�d<�\y� `%�N�;�W���L~���V�����!÷��h8���C���$3J@+)�&d�����6쟸�|b�x/�[�_�N-�ir����5(H6�3�jP�[)��m�l+��:�t+5u�;(�f#���e��t�PHM �J�p����#
Z��t�L9��6$�)��mC琡��+6d�0K�g'	���r��	��H��ݤ����Co�V���1�ʥ��@��� ��Y�'��i�����e5~�xP�ݩ��K��fD���a��0Y�?tU�~|9�1�����\�Ȇ֔ճ�,c^	L�$�F�x7�&��<~�l�3�r�2�0�����A��1'
��g0Ҟ�������}�-T�ƣ�S�zź���}��84?ϖ;>�:'�ܷ~w���q�`�y��`�E"*if��X��{2�p?��RCB��2��&eW�ö R��Q��Z�	"�̒!��4j�>6���d[�lp��^
Ys�E3��d��_�R}���bk��XKa�tǮ\�~�>�~��#e�L���@'�Q2c�5G��e6]{9��@ּ��s$��{w�����B�v��g7�U�;�����d��Dd�K��m�h�^�הPǱ�y�4A�Rn�򶼴{l�4*b��%\T����nؔ볥Dw�ʃx#
yh�/h��.G���?I��,���]�s��bu���(߇�V �k����p䦀���� }�N&e	�W���)�5Є���,(ܕ外�0>��N�\��.��?r��c�:�Qq��Drm���S�8Km��,��B-�'m�m�>�<�#Jj��W�}r��)*bˊ�W�1oŚN1b^�1���)U�X��: �]/�, ����]�HO��3��J� 1A6<4)��p���
�����#=��^��&���%P�oC����^��EA䌨r�;o1�� �����A�@ʛ�24R��F=��MY�fc���V�a���δ�U�eia��
�y��i�߳�S	��3و}��r�'\� �ApN86H	��?؏��Ԙ=vB"T�!v�vE7��A%�3n򵮸V:ܑ��jN�g'�"J8�x����sG[�YӹD*��n%���@Nm]�Z��x�6e�moi�u�yR�o���Nem3�6*�����#�ŷ�Kɜ3
���1�t����A��3~�&�p��#�B�EUH9����ǘzI�U�S0Vn��0�=���ւSo�U��!�s�笗�Ig!��/�l���)����A��
�*`"�i����!�ܧ��@�MW����1�����J��d�z�aH>�+�A8׈��<t��ഄA��y���2�2H���>��>��@�g�S�P��=TOA�:Wޛ�.L�r��n��������D��W�nx$��<<��x�����8�U��H(�{�?����� ����}_R�D�%���퐳V֜���5�i�t@&}�E�f<��Y���ۻ�ϱ��?�ku|�8)�Z��{<𩀸�iN(�O�q��ܯ&����¸�K��c�w>̾h\�����JA�y��!ko8P�{�5���^��f �����׮��I���q��5�q�0~�>���Q��L��:'ԙ-%$k���JL�Ng}q�Y��p�4}��o��3��(�׍�o�2.���C���A��S'��uk<��c�2���O� dMU�s�m3 mH��<� �� ��ƃY+���n�聅��a��W5�u��\�i��a�%nI�f��s{��K� ����\Z��a��i9-�n�����6�]�x(�}A�*���:0@�6���<�A��"�
(���ޓ��BMF+�l���qC�-1[�.5����SZ��x�/z���)��w��OQ�� �*> �+X�)�-��e�q0�9� �O!=��|���/y�_m��S q��rW`�^������XX$	V,#��b9�| ���1�-��ɄW�sě�����@8�`��Ә