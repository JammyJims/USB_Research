XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��=8u>LG��ip��f����h��@p"����(�i�)P�̲��T�\���	�A�g���NlV�Вr~.^�@l��1�/\������[Γj�(`o��a���"���>�,��@�����Zn�{�i(�.���f����?Wkv����v�>��t�[��P�|��-0������3���&�W��E�6χ�O�"�.���nvˏp?��߅z�c7��9R��
�H�4�q�����֫�����fw_�8�U���Z��t[tR�{zoak��6�ߴ]V�Q6$t��b��ݧ���g���VAg�2�8��c[��n�a����oٔf.��N��I+�ږ�e%���cZ]�j0��!`B#���U팍�u���	�3��\�4U��qt��&w�8�N"�	��W��.��,hF���2��BV`Yп)}D�N����M�{�P������J=��f8<�C?��o����kYk�>��t�3Vj�|����-ފ�P<o����E����>w�ʙ;ɹ��顁�m4鲍繘1�� U���G^��0J��q�ս0���`��Gw�Z߬�cO�]�O"�$�`�����*�z���N��xM��.c�R!y�'��?�o�m]�;��I�{E��Լ>J9�6�������J���g���� �q���WJ���ߏh����1N!2�  @l,l�^G�����m��t:���{*���|-�g�Lr3�����SW����MCa�dȐ��M��9�&�VPZ�XlxVHYEB    2a84     ec0s>r��掰_ .��,.�7���Y״΄5o���4�{d�1+���^�P[�=kb��&G,�'��܏w���T�	�#�>��
�"�=���aSlO��D;��楼�6Iq�D�Tz|�b-�Y�H��"B\�Y��L}� m�|ų �Qz"��A�4jQu
��a����o�s��Q*�@�:���Qaْ��J:�D-ψ Ŕ��F�(F2�l u���R��!����=&�9m�w��;�0+�6a��607��F�Pj���WI�8��{�Z$�)�^"�I�t�*ʩ��q6��b�G񱵌s|0Q\�CK��_�^�=�ĥ�SRi}�Q��lb�L��<o\4}��=O���}8��d��60c���r"���<m��b�3&Q��R�IA��D�E��*5ؖ��S�hIN w|*5ɮ6��s ^@���[�f�t�'2g�����|���tVpM�[
�*��q�ѪN����*�0,�OS���FZ���rn�d���|�(:-Ҥ?�I�'���u���>�{���[w$S8�ȉ�m��ٺ��vCY���w�N�PL�ѮW#����U�kGӨ̏��t�(F'GX�� �0}�N1�|`Н�������8q���|B�}���}<o�Y��D���8�+��[��벒!"]��R|xv5d\��x�r�9W�>��o$�emYy����H��S��=1�6>P �BRm�MH"��)�����ԕ�D*�]���Ș��K@�΢�d��X�W�يgLq ��@ajXPB�m�E;���X��*�Y����Ly�����<Nu��c<��n�9p�p��zm�|�R��}�Gq����I|��	�y���K����I�i��_ //!��c!�'#����5�f�����}��cfV����V��T��2X�z�,�B���	%�=�"ӛ�	�Zu���@�iw�f1�'����S�FjW���v�˙&G7n fK�]Y♢��DۣA�������>^d˅��x`�mfW���7��]��Χ�g0š.�n�����vٝae�/�l�wq��P�W"{��Q-ϭ�2���B�v��FB(&��W�`)��[��M��8�Sġ��oX��7�6�����B�pr�$���ɟvy�]5	g����%so����������~(��m����+�)"vj��0���i�nn�y�Sjx����A�b��j�� B�[9]&��Q������ڕK��򯀡?\��X�_(��,)��U��E3���&6{��/�Jś
��ˌ|�44�� C9'�IǇp�=Lc�>z�veI���FIr?^o#���ü�}�<��׏�m?��$�T�L�L��1.�������)W��e���h�I_���	.�>�X0�וD��l7�`�>��f�`V@j���~ �����ދ�l�=F���u�Iýc	'6�&�՚��q	���D���Er��@���dA# m���u�`QH��`$>��7��Ǎ�������G["�|����Qi�b2]��8�,@��3�Cq��t�x�q*�3%I�n+��ڦ���
������K��X�˻CZvI<X�d&�CI�'��I��Z�w����l�R�r��w�-�4����'zޏ'Գ��.uk+�
��L��1>j�;��=�k�y]�C]�	Q
¼f��L�LGr̮'��O����&���5(�����6���۶!�I!*��q-L�dj��R߮��HV�(��n̮��Ԧ�� 9���zI��\�Yj8l*Y>�a%�]k�?�)��9Mlf��
���n����$�B����Tw�iV���~��4�� ��0��9��`w����	����+zC�b��?(2z^Ou~D���1M�:�|i���Bl,��潍�D��HoʶBEh6��?�XU��縭0�cJ�+l��9w9]L��^l��H���ɔ{�Pu��M9���,��H�i��;��k^�4�}��!��=e%����"�{��jn�v�d��3�9ц��/ ���^�aY���B�j� ��o�A��l�>*LC����Ү�n�kÕЭ�^�E��M�č5�,S3���\^��
��0έF��Y�1���ʈoS,���,|��'�D6Hw�^���z��a�����^Ds�Ӫ�iK?��tmL�_?�q�Sފp^rA��;��ckW�����JrOQOXL�|Y�����F�A��U	���lͤz�KTD$,���_�a+w�L��w�d�� ����F��/!���)Ҿ'_B�y����+�|��\TJ�*HB;��m@�����1��Y���t3r�z.���D�낞.
5���3�iJ�s�F�H��}�:��r�eۺ�	:7 ӟ͇��6]^��&7�2!3�}�5M4�s��?�H�� ��׭�Qt�Ƃٛ�@��ǟ��K�_���@��̬��]��/�8�wz�(�b-��rX`n.��L����������u+u,������G��L$��\�w�,���T>-f�tG3���euwK�U�r�7�eC���:���&�)(��U�=���Ԛ�&c�f�$�����VƮ]]&;nS�|Gy�M�<΁5�Z�E<0�H ��K/1��k|OGQ@kWg���QN�J$�?}g����qtr|C�w?<-�1��\wH�*`4�:YU/tI���hɅ!��&X���-�t��1�Gؑ%�n�}#9��dev��x�  M9R�Yr��r��` 𾲯�DW�CJ$Uv����j��%�h���^
�.�Ҩ�F��d��X*�%�"����X�R���'wp�r����S`5�F��L�`�R�°7ef�
^�P��9���P4�R�P�Z��!��}��~���Q�`�nʫ<vU�L��x�cve���x�9?��y������k�X��aP��]a̰�S��J5���bt{���l?/~������ˣ
-?�'3n;4����8����{���� w-է�梨��(u��ʦ	�� ��wq��x��ί���9| ����B
�X���0L�fxF7�(U_��N�����Y�_5�ȎM>� ����%ɬ2r`܉��ӆ�@Ȇ\��J�L ��2U��4��S�f���%"���A�J{Bn����2�3�c�0@���S 1k��Tr���=ޮ���w�Cc���X��"O�P�g(��7v}�{��yAX�rE�C�C0���e@�;5��>ft��{r<�;���;w_��!v���W�
�C�%��(?��
�����ؕ�;�A��D�X�6`N����� Z�Q=�2�v�^:vqוD�˅�um�U9��Tb
�GQQ����qy;j	c�{r-�ff�g�/\�J�`�����*�9F��������ʥ�u	�ԑ9<�&y��UzgX���U�[�o&|��\{z{9�Q��K�����Z#(;iw_ӒZ��E��ܥ9u@�� ��	���ф��[�A�b��4w&�bt�I1껩�v��B}��SpҒ�������:��2%MX�.�?����<��}�q,r��!�cs�&
���S$s�t3���Y�^�"<_.$�q��>s�T�ç��_�봹��}iğ�DF�߭ݓO����<S�D9�ĭ�um�C�31%�%�eP�&`F�b�!��x�:5�q9�"X6`�����T� X*v,^:q�����������Na���