XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ڶ�"t[
1�����';�*�V�̙"0��^,O��,�H��J�G0���D��������S�b����"���ڶ�ɄH��`��ޥO7k��tS�_3Wd�Kʂ���P�O�@]5]� ���y�d���܃���KˡA	3��VV�7�r9B�s�z��7��E�;e&�3w��
�Eǉ�.ϋ�@���pD���XI$7$����y#~��]TT`sbZ�SQ������&�٧P�i�����=�Z��k2�0(�>iaޥ"�'��|÷��^z����k �1d��;槣o�d���J��r�$/�Ϋ�^ $��1ZI�8y T�^���#Q�U���g�f����vcq�4��k���@\���%�>�I�B��dG��Oѫ:Α�aS�Xf2]>�eö�J�c`#|����+Bo���m	�U�0�
�����b�Sq�_:�c����)�#_�!'R�'�ԦZ�E;��hKB��	��O��{�k�Ý��kH���}�C����Vh}�9����p��$+7�6!V/�
y��u��/��鋓�[r5�Ʊܭ�R6"n5O^���	s��j'��-�c�n��)�� �H�en.��*\x���\ y]B
���j5����%������y��g�:w�$�����Xz5d�('�>X&9�7<ь����,:+�t���Q���Ni^q���Sng�5S�oΨ�P��G�HC�( ��؁ pb:���N�=־vQaJ�#@X	z��ت�j2XlxVHYEB    2901     af0�#���=؁^*�v��?�Ao��7��ܲt�c=Ɂ�Z"'�}�t�Ѭ"s�-`��yPy��n,~�f��HQeƑ�Rblru��;�=��A��)J��y(-]M��i *2J�p*r������(a$4�R�/����~�0�!�L�_�{��)�A��l�A�/���{��V���æɅ<^�:o*2Ҝݙ�1z����f���RZ\��𼟊��R1���P���&oaLxQ��c(m�d`�l(����\�M�T���N����G��[j�����Q��Y��/��� �v�Zff
�!vF���gh@lk�L�����&������bߐ����Д�,�S��?�	Ǿ&��J���['�����@Hg����le���\˚n	Xn��6+�j��n���
�.����a����O�w˱M���Bӄ�����o�m����{u)�Ѿ�@�V3�k%+�_��EËe��� �KY���,j��e��G� �8����E�uZ�Z ��b�&����Q&!��:DوSI���ڴ�`���5V����8R�D����dx��E�^��C\7�}�:���e�j<'�%�,�]��pl���.��Z�h�C�TS��e$7J�m�A�`�Z�b���/� Olu��<9ݜ&O}�5DW�L>�vEU�qT�0d��n�G|����t˷�h-��b��t�;�-Z�ԍs
 �^@1~[Fݩj�M�6��.��^�z�P iVX1X->����T=?�P1<y����~����C�bls��b8�Q˓����t�btT�	Xk�����`&����Q�3XY�0�U�E��o����at}��ҩ2���xK�خN;N��?iԨ}�oqO�X�e�X���5��+� w"�b�_@��C�ҕ��ҙ��5j��-�+�ˊ�_��+ԟ�r��b0���.:a��E�t��	@�C��j��ʗY�z1��q0�d|Ih7��-
��?�aH��=�&|�d�M�OP�i�P�o���.�ȸp}�!� ��y����\~��E�Q(Vq��	��q_�bK����L��i'/K`��oX=H�\a������ףX��+ө�����{h�Ѥ]T�~f�C��]%��	�S�+�dr�Rh=��a�ZA`^,��RU��V,s56WUgdF��<Q��p2�\K_#|���9̱z:;�m&(> 4�$}S��'Jm�hM]n�n��V��L�:4ӎ�O�D�4Jsao1]�F�=\�h�6�	��4�x�V0� �iʽ�}�ۻ��tx� $u,z;��Z�� ��~�(J@�5�CZ�Iht�ׄ��EyB��]�M7"��!�U���6���%M3M(�̥��nsXWo� ����A�YI��j�ՁT��-��vR����׳���A�4ɳ��dJ1<p��=��o�ot:_��%
>�g��Cv�4�Xο}I�3��-�K\|���7譇 AݽT8%3���X�v(���~����2iL�ي�-�$��c|E����@���݃�����e��x�~�I�{��N���v����0���z���-x�j�K,�#�QRm��	됞qX&������
��]}O;k���o�l�~��'�$lt!���Q�\h}�gG�������PٔkE��"�O�� G�UG�ַ��ف�ԫ�[Pg��C\zeCl���ŧ2��z�To�i�c�u��� ٠B�n�F;�3�NPA	�)�Xc�AZKT�}��8dWJ�.jt6��U����
��/�5�'	%�|�u
���L��Q�	��9�mb�j����H����SF.Ę��x���
['��Lc0n-�c�L9 �#�����H�Qu�����[�|"�s����h2Ļ=G������,<���}o�$��po	2U�}]�� �D�b}�s�]K��:%@~����
,��͸��[�s��s�O��eV% ��$Pdt�ɧmyW<�� ׸�'��8���:�BK��Ԭ��lP��$���&�^�G���v�I�W&����%����#ޠ�0a�&*O*�K&-$u��qm'������^/n ߃��A�~I��+���G��%���.�Ne�>=��~�0��&��}8�G���!�t�3	��o-�~Sk�!�/��Yg��~�h�&$p�&t�%l
��h3(������v�e����t�.$=m�yK�\�߹�1%C$Vy�p*�.������S+���ɫ^춻5;kY�IPNs�lW��%<ۛK�Ư+[b.�	��"�s���.�I�V�(��{�_n��$7j���㻖�`�ǀ�U�Q�.�$V�|������#PS[�m�DЍ�a<��v��2͛��7l��%8~��hʊV�ـy�a��ZKt�7��Xǈ@<�p��6|�?L*k�f��3�~a�2��R�pX���<>�L��	U���+�D���@�9�ޅ�j�q�v��(b�����|<PM_$��}��8v�S"�o��$&���
����M��[]#4�<b)��(G��	�ǭ�C։��2p]y�ʽ?��]48�`�� �q�������0?~?�%�0]�#'��6W}6{��U\�Һ0=%�>��w���8Q���Ƅ���n��8(��Kb�e��q��H2}M1�M�X�PEJ�*��47�����a���s�g����f��0G�Y�b�m!o��_�Q��B�M�"t�\U����Gh��BaZc_��ߚB��äu�7�b����FB�J��V�t'/f�%���6���5