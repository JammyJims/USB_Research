XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>���=K�
���)TE+�#3�p
��[�,{S՝Uu����C3s�.uS,(o,��i����&�^5�>u�d�e��'��ƥ��[�z@��[i� �z��#�x���͊�Q�����ۛ����� ,e��tŲ�.7�s�{��Fۏ({N�^^����$M��3Z�(�;*ݶ��p�_>�V�� ���0����'C7w{4�O�w9<�7޽�>�f��t�7e`��b�m��H�	\���R�hj|*��Ѭ<K5n�v�_��4���PU<��&M}���J��o�œ�`�w�0�Q�h{Y�˜�����97��U=����
KoJ���d[�]O67Vu��/���J�g ��}�&���Z $L�˂�>�A���S�{�q+��77�5�j*�Ώ!�wSt�E&C�-�J��2�q$�?A�l��t��P
'���~Z| �2�Eԁ>"" =��<�N �ߩ�/�On�b#�� .u�l�o�9E�W1����?k��6�|
�+���ó�ֱ�V��iU%�}w]%�$`��EM�=�sZ!j��*���eʩ�3�E�jbBMW	��G����rzm�D�����d3f��k*����;���H�,%�Ι'"A���Q*	O[�?׶����BE�����[|�K��|zP�w�:��W`�{tOӚ݁؞�C�����oq��>�����iW`���[.���Q,:�r�h9�7'к��� ��ާJ{���*y��ڈ�t��v�XlxVHYEB    1dce     b50L+ݻ;��_��͸�b�jd���(D�{'إ�gR�w	�{R']�P-��$&Rb\`���_�Ct�fE9Y�>y�P�V�JO DP�&f9Z������R�����L�L)c	���WG��A�D,��9��}���?^.��Y�kg)�V�6�r�ʉ����r��[sm9�z
]w�l�n�V/ھLQe6��5�鞀�9L<y�o�c��QY��Y稖%(`zN�U��4���"RH��[&�n���ݦp��FGN
��?0�$�u�D��7E�%Z٬�o��rP,='��+�rg��}�Dk��z�
mDq�CuNL����2�!9e�a�M(�Fw_�&��-l���rH��Y���7���E$�[���Ҙ���]&W�e�����L,�$�8��3����4˲6�#�z���!�<T�'&���&��.�_�&��k1Ae�Ş��܍;�
%�i���͔#D��:J��0�ݍ�c��/XIII��Kƪ����II+Vۙ��F2��8���;�\V����n��9���LU`+��z�Эg�Q��FL'��-x��gT~��4�U������s��E��ۤ1P7�b�d�8П��J8l�����_��ͬ��A�6�D �þX<�)f.wt*�����I�+��Ѫ�Qﲎٗ�4m
SI�5�(�>�!�˨@�fm�g���r��$�b0`��<p<#�����HOJ��?oG{�����-�P,��ڎ~i�����Q7���s�I�E1�!�*�F��QA�5�/orY	#������
�����!�q��g����f�@ VǄ�f�3.�5A)�Ie{��}Xk$�a��!O��uE����*��[��Y���9�֫��qwV�[Пp#���Qx!k����T�9A�t�,0듟��WhE�7�4X�o�Q��!F�����z�!8o�J�Y����Ԓ�t��6fqJv������d�08<��Ԙ��]�nKy��ғ�r7,�lY�!�1��rʍ�_�=ۤ;5�N�+�.�v7uI\+�t�z�ڄtCc��2 �����F�w���hQ�������E�o�GL;��%Wr1�~�W��� �yD��;���r�zP: �?������3�I�9���(.#K�M�դ7�����A��裬��M
�D�TYdgd�=Q+������rv�[��ST�h�z�쬑����̐}G�X�N��xN2��y�
Ooüӟ�c�����[���}�z��a��ʽ%@�&���P7���\nS+pC�H�s�6��cB�tc7U���� �	�ǪB���L�$��0�_��������	/��\c]���=$��w���e�&��,Io&� O�r��2�N�&&���;��hP�+���Ac)�x�?^�����>$i�� �ҟ�!��2��Ai�6T���X������=�YFU��Ľ�n��W�����s��0r�BɅy
}�D�␺t���twFr��e
��Zl�:z�f��NBEy�ˮ?��΂�S���s1�}�}�J�a��U���',�
ծUmp2�}�vA�"I��EOǗ���e�/�JL0�j<�y�D%���S���y�����W@1顀�w=O{�?��u`�9� [2X�B���n#�����D3dq���Q��y�>�v|���_����E7|�#���y�F�ɉ��K:s�r��_[��+��4��&�5\%1	«�����p�L�������:�Z�ɫ��;E�["�����k�ې���e��{�"'�1��6�Nr��\���Ʀ�l9@��Ԟb}m@}�T"JuI��q h�7ѫs�řW��濫�Z�?6_Z7�T�
ѻ�څ�'(3%�~ 7�QS��&�W\ZPy�'�i���������J�܈t)��������=zL��qiK��g�Pbm֘E��i����\��d�m2ߐj|t[�F%d͑��O����0���%�F��b��~kZ�:�r	P�t1�l���A�}��� `���M��7R�VF�t6Z�����eR��ͥѿ�������
S���1{N��I��=S��=0��##~�F�Q�U���$�w���S�Lv� x�2��-���� �|x� �cw�Z�1nD}�P9�C���C���2n�SJ#) �\�^ө1$��/4g@E �p	T�f{@g�ӄ�ݨ�֐@����,_O�O=Ǭ�.�O����RGtd���e}�_斛]���v{�d�����m�;���x���z�f�͵ ��aZñ�)�5�!<4���_��__�&��{���F��齸/ݑ��]��Z�YZ��[떎߬�� ��4�P!�_|dV,��2P�vs���6寂��p6��j��f^�3M`4H������������,z�O�B�	��"A�g�{���K*޳p�f�ӛt"uh���j!u߱���h�.��i���	/��9��K���0��H���/<�a���A�� ��03M��0�������tg�Ւ�kʮ�'��  �Њ6��h�/A����"?�qy�O�Y\��=���Y�0�-��tDw���Fؒ�)��9�H
d���	�+��Wr�*�Cu���<QYc'zy ؃�J�_�ð���I�H�J��Q���.f��ݙӛô����g)�T�/^l@����:�V#n	����Քjm�Oƾ�W*��`�4��qo����r���|'i��z�c��ya$�ӠuV+EVW���P�2���D2��S�2����<�/$5ǎL��
�6�Z�$�O��;�]Z�Ġ����-t�l�?#���t�]��T�
�j�+��o���$GLi�����'J�/鱟��{V�XjG��4�