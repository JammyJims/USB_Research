XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��IO��xU�DG�[ſzu��H6��V���/���,���R�v	�^���b�,2����)0fЛN#ߠ��d^�ū�!�q�{~��Ҝ���"�F�+feʵz�A�`�'��_�7CV�a�����j��5�IU}��8|�aʆ�F+���.6��<�U-Ɏ����c�{�����É�P�8@��v������R��j��L���I���Z��tef��F;�0+�٫)Z�y�\�b#�R�Y Ȍ.�5{����/j�����a�J�O���p�4}�3a&$���{���j��W��m�1���DIe���k���x%��:F�l�ʾI�ΚT�m�|�N�����j�3]�j�,�p�}�&'t�� �n:��$����]c	���Y��ۖ�d*�u�K���J��BهZʌ.�Q��n�8��V�8_�tX�q����vM���|�UP9���S%�4�_Ş5�	��}����/��'�:�n��4��i��Z����|6��Gب�E'��B��c�.>�2�E���	���#둩�:N�c��v D�ר~�,�(�2?�f`7��&��i�ñl�5�g�G"������=��� ~��`�+�xX�������'J2.�~���4�|;��bZ���#pv����T��~�B_���Xuk7�CνD7 ���c(�Sw���]I�`��9��d��y�a�T�`s�Dp�����$�ı���H+|�C	3�SQV��q��`>���XlxVHYEB    1b98     990ǥ?���6��g�ߦ�k���[�T]Rg��1���k���^~���k<�{IC*���(��IgEy��WV`�������ʵ�	a�3W/�r&:%m�<��GO޳m����N���U��jHr��a��Z�`��� �W�#�Xݻ�����ˉ����+�+XB1Ӊ��t����^7�f{&"��\t��p�	��!Gr-�$�/>���ځ��'%���Q�����ݓ
�3�9i4�=����LӔ�˳����.����N_��g�k�� ߊ�:]����d����/��\Yy�(�|TW��7��y�/O��5g|�������t�Pc)N��ɬ˿/��*�F���8��Aۏ�Z�X�.:�ʘ����g��]��vS�i��o�pPV���
����JA>��� �N?��i�%��]��x�vJ�	���~��6�
�������v6q���н��I�!�0*C�����z��*�RK�ŕ}ہ=i*[x;���Aw(�6=x�]9ܛ���A7c߃��m嬤^�^COJ�_XN�+��Hл>�J��Hz����.�)+�_���*Z�Q!�]��43=I��_��{A���8�T{�Q�mZ��2;b�d2��@�{�m���!5t\�ĥ��$ ]Ck�]���D��/c�������ü�9�D8����7�A�42�6TCD��ӓ2
�P�ʌF�փ'�v�[��2��D�����"_�������?A=ako�kI��#�^Q)�'�ד�Il�{���E?��)�z��`o���N�5v��P�f���k�ͯ)���B� �Nt���
5R�2}���%{��Q�z4UQ��Z�Ϫ!$r4�.W��&����x{�<��^*7]-��jL���<t�ےJ\�R=��ֺ1|��K	��[+3>zK`�+ �[���L���ן��^Ϟ�A�I�U���J�h�
`�R/z�k^���¥٬�-',�T�ŉh�����|��6-?-��y�n��*s�]�q lNr���+'}(� &�F[I|p�2Q�xE�~*'�K"�T໻H\(KژG�W"NP?]%�u��[N����E{S
Ww�+�]C���,�dS�j�:����^0�ߨ,T[�t��ҩ�� �A-S^Y�Չ��Q�w "�p�42vvD[aW	Á��74;����s�F�tiXD�2�a�wfj��J�w�7�t����N��F���EP���A���-Ch���3��\�0�s��˔|�B#ڣ�Ti�,<�[i9���+_�Gbm�Tbd�|澈�[�&ܮ.I���_@ �1�.}��� ��G��?�W��K�K=&��Q�����AU�)ESq��A��u��8�ZG��+KPЕ��K*�ĸJ\�����޺�R�!�<����D�w�uC_X�����\��;��"�^I�t�뗶i����b}��V���/�^h����+ܬk\@���:��69��#@��9X��+��E��:+Ƴ\��b�[����zo�'�Ở{��x+�A���pJe��5����:Kn�'����y�*Fl>��������"|~ݬ,>�&��I��"%���� >�M{-E�Z��~	o7
�{�u���*��0��@��c��BQa�G���3S[�2�ϖu�u'o.v�9��pح$S�-��xb��[����S�+��(�[�<���9]da(����fk����1���
x�.+�f|{d��;�dT��F�2��#��������DȞ-��}��^I�¶�UaZ�=yW��"e���*�/f�ӑ��z�|d�UuȠz����B��W�<U�L�:�e3�c�	#nƕ��2
�xO�-����uO
3���#��Pds�ǱA��'H�#�I��H��N�!+�39����p��j��A �dۙ���;��)H�޿B�&)��؅�S��ȵ�Ѕp=�_�uj��`R�����3q�S��~�j��DN��:��s!�-Q$�����!�CC����������T�6�*9ݬ����й��t5b�$g�7��SX���TT��N�ih_�J�R��~� ���Բ���o�v�/����e}���0� �~����,%�w�G�g�K$��?��U��t�>�<b7^�Y:��Q5$f�6�F�ۢ�.馰ޏ��"����Ub�=
�f�9fHU�ݾ���F�����_� �O���U܉�ăTRh�}��3H�'��Ɉ�NC�B��~�X�r�C�+X�(J��a}�<��;���T8s	�EUT<�w�PKs�=$[������1���YG�:8�Z��,��"SD<˩�$(0����f��\�a\��_�n`Y��-���ߑD��ҙ@��1sDt~��H%�y�q8j����2�AVSz�T�% bpOWH���V\r+ͼ���C��B