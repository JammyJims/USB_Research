XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�"s���Ŏ0�ŷ/�Ɯ�,�զ���RGN�5��v��ǫ~�pV�C�K�3����؏�O(�L ��8�e�O��ݶ�%�o�o�����m��a���h̏�G��\)P���Lo�]�ūK�̒$@I%*��I���_kT�Y 6��_�����1�H�.W0�:=��բ������ɂ�/�:4��:�w�c>�e:;�"q�$ٖ���#���s!�p�b�r� �V�ۣV*M�}#R��c �d�ŵ��
¢LH\�G��-݀q+�`+�-�1�oI�*����{�4Ӈ�7�F�G����mU���"9R��^u�7�L&-B��BL ������}����0Ε���_��F�p����@g�B�ʸ2h�a���kـ8|R34N
����'�m��<(�N��&E��čՀ���uJ�=0�VF� C�ޚ$�ˀ'�I�h�q���3�7)x�)��<�V�L�m���	v�n)3�`��ע���z���N��%�u�m���[��<��0��g5�p~��`�������W�piZ��=m 쐟�]0����`ǖԊ��ї�{��ڴ�ߟ�{m�څV.d���d�B7�.�y������Y<K����Uӳ�}� �����K��Z`�]ņ(��!jbܣc�T���2۸ٯ�VT����U$ڰzt���D+�b�����ų�T�iW'hpI�d�N���ɯ�8A�:_GH�xz0��h�`o� �
_4�9ބ������W���z�
��R1�S���XlxVHYEB    1543     750��k�g,XΌ�֯���a��ڧ�pA��~���z �2 y�z^�r����:�po���)�P�A?ΓK�A�u�"J�q���P�b���Fg%ֱ���u���v�����S{�E�ĳ5NդI��B3�eޓ*�Ւρջg�f�̌���S�z~�ݢk�ۣ�����Qx��!ǩҦ�]�6��V��[C(4�PȾ��GOiȊ���vݼƘ�1.�H����U�s��J� `3�r2+/M���A
�,7>L�<y�f��SBS(
?[��5���9_o:4��p�=��6ª��tjK���*/P��5R&���ﴱ՛�a��vh4�X��i���D��)���D��	Y ��N�_�l����� ���=�C6�*e�7f�X)T���U#�0������

4s	n����gRV)n_B�����kO�UɦC���uiXH��4(��N1Q3�]Bc�3�i/讎$ �.��v
S���(�4sfZ ����c��(��f���as���p=1^,�Ku�B ��4�p�;�a,%U9I}L^J��J6�E6C�b����2N��ލ�<n���٣ڲK���#p�u��s�k�Iq$ �w���9����+
̪\ �ׁM0�e�Bm�A�j������f�*�c��n▰��B���_��4S4����F��=�V�98�N�l��ȯ{nibO��}�~��RK3��s����ˉמ���N��=������ՠ�����eS֞�@'�Ί�`LUx]%���o���FTV{L~$�*����&��N�,�UK�(=��vw.:��o[Y84߉����`�K��gas[O���V���44(�*Y��؇���s�nf�1�5�z�/�.=y�7��
�x�1�9"Vz2 �&h[��G�Z���C̎Ud��P�;��Pi���tMx܁4&����+Y�����ţ�x��(|T �C�f�)cq9���I�u�Bs��]>�в��~����jR�~�-�!���G�_���&#��J����4ٱa/yW�+p%{�&��TqQ3�{������Ӳ�6�Z�}c8W�x��W ^��h76�A8,��k��]̰��CW�S皡vw�� �����XV��O��4�^��|c�@Q�8#VȠ�=-h�� �'�� m��-uN�;��)�������[�Y�K@���zm�[js����uRo�$�υ$H�=|skd�3&r
mC'ꤨ�K�1K_1�[ak�@������%�����Y��Q8���,0��%���fpu˥!�͠�9)����ې&�(f��)W������?em�����v�6��h1o�Dr����s�EpPbޖ�_
$Uy,"���'�X�x1CDWe�σ�no�V�.�3����D�A]�Zk�ʥ��s?�ɠN���B�=�b� 3�bS=m�\Y���Cu�=����E,��K3	|�S��3�˩�a;;}56u�>�;C��-L�����;T���V�E����h��wJv4Tz�Be�]��+�tPJ������Ti�E+����s�T��ņ��g��+��f/�Tg:,o�M�3��j�QDB�,������Ӱ�}OGO�:EܕN��=����+����a�$ħ4bu؁�������)�]��C�m�����r(�r܃�^r��"�)�{wP��<3�����T0Y�y��U% E>\�f�:�or�[3��z��Q���� t�Y��zbR���z��F�B�Xq�-<(�	_��z'y���n��zU_�O�X��'���D˭�.ڏ��}�y�ἣIf���Sl���bbfX�Ng�yU̸�= �B��4r;��;Ï���r���
-�hX����