XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l�����e���A�f]���MkF����w�H�����p����d�������D��\��ҵV����h};L���a��g(� d��:�$J���9}޶]��bB����?���d־Uy��P���\B�S��2(�w�Ƨ�F�>М����#�I��*DX�V�>v��� B[���/;M:=L:;����v:�i����M��0\�܇�$ߞv�)�2�\�ɢ��r��w୑%��7�GvEm͌��>�y�:oY�h�Af}5U�M�o���!��}���M?!Oվ�u�hy[#	>�P:�P�T�_���")I惉���]z��t�ET)FM@w����5��݈�0�bצ+�2�P,q���b�ZdO+ř>'Q���D`��	J������?�3�R�tZ�1�K(������GX�Y3=i�־-a���l*O�q�y"�-B瞞G����g����%��<�Vq׫d�v_�:Dԁ��лwNd<L"�c��n	5s ��-�{�|�2�͈*|���x�Na!l��fVP���k��籅�`�Bs;�h��7�;�/h��q�=n$������m���r�W�獳�u5h�V��ǒ�"��W���l	L{���Z�f���T��H�|��*Ȟ�}�·bi�IJdA:��5Hqf+�o�w �U�ַ��V�٘��څэ�J6�Z��mh�	G�ՏP���?D�����+7N��#@Fq���yN�ŉ�~U�1�ȶ?�F���r��'h�?{GHXlxVHYEB    3b1e     db0��_����Ь�z�"�����`�ș�)��o�"���6��QW����&����_���.��,.��0#Ĥ�$��ܭ����c��6���nQ?i�z�DT[Yw����K� Z���P�sS R1$I�B��	~]�Nr�J��F{Fv��i�����r�x�}�a]�d��٨�N�"�	*;K����� ��p��;R��`��ո4G�``ܛ
��-�N8���;"�l%�M����b�P�(o��^�ꚧ8��U(� �5k~�r=��]�S�.�^�=���^�7p��$�2�"Ud޳�d 
��H-�M�b��I\^����_��Dp��#T'��;���Lq ǥ��[݈����0M�WF`��%s�q֗�y ';�L�Z���\㲃���~oV�Tɀ����4�fD���N0�O9��w��*7�@Y�4��su4��S p��S9���]��5�OW�ZF~C�A�zl��?�!x/w�ۍ�$�>�q�R���Ta�a�,}n�i�3�@�U��j,T�I�+��7@aĝ75m`���/?�=9N�E8�I|�J��G=�����=���|fVn��	�Za����1R��rr>p'GM�wB���PB�4,�����SCw��4�[�o�;uE�1��@W�eis.�0��}��1�7B�B'�݈�s�p�웜�2��yuq5�"0����s�'yM$\6!�cUq8�|���gy˽�Q��\	�
ҫxGF��6�`���˃j'��=�#�q���3�m���u��C�H���������?�%XX���Xe9�n;��V0�A-��[1�LR�Գe�]��ȵ��^d�U��~x"�TS�:CС��v	5���$� �<]� B��;kz��>_{�8Ǚ\��@��$�U�͘3q�����n��n�C�/5d�vHMʴF����`���A x���P]�OLg�s�F��O�?�Rƹ��H\�@ܐw>��Y
�ms�:I/�����Ui���~��q�Ѹ�jY͌�QXka���RՓ��s#mb�x^���|1m���Y�ƛ��Y>^�(�9�[&�yaB˾q�KmV���������i, rzUo��脾g���ǔYKq^`[��}c*�,��#���x��Ⱥ�:eBm>FOǷ�43˶��w��Ϯ�;��9�?v�PY�Pf.�$��0���y���W�Zr���W��!:�5�s��s�գ�l��:ؠ� ��ARO�ӈ�ޡl:��'l���&�m^�ʜ�j4�Ծ��ݼа�睼{s�2~m��.���k�����t�B�5�Gs��M�Y�:���ym-��	����%˨�i.�B�j�u�W&sYޠ)Kr;R��-5	8�O�p�=`�s���-!��Q+߿PQ5���p邉��=���(�{v��B� X.�W���?��Gt�ٌl��8�.�{�	���'�8��Ј����D�Z�Y=����3�6�
b X��F��BSWĀ��z�n�[c�ϝ1�`,l}'��f��Z!�I]e����x�j���MيS�[ ������C-C"�pR5W�n<��6+���ap���~�3�.��v^��(�k
���k����wV�ǒ?�r�#.���(��ĝU&Ѹ�yC�R�G:�n+�<}�c���;�5�))�%�_ 3Z��G֗c�^�X��?���I�W�-�z����DAp�� �(�Q߀c��8;#��6t�g���j��[�p��Xj�
E�L4F�D��Sb�J��� T��]
�:M�ک^�@w��C>�4[a���Ly��@�+�:Li�F��1S� �]�I%�y���U��84�:#x��rf���1lEk�0�-
�3@��	��� �6���qiBc�U_l���g�*�2oM˩��bo��YC��S���ߧ�w�17TUrz�S��Ok̘X��#��)�Y�X�$��X�5"${�G_�/�Aa������f���d���)�W���`�M�\:�j������\(�9�o��q1�ڄ�V���֭��$$<���A�/���z�͛E�V|��o���`�p2}��W��-e����W ����``�����"LN8�@�N�1�S�(��S>�k)�d���m�sKq�	�?� Q��ob�g�����A��*bVEח�v�K�`0������r	�+zc��o�ٛ��[����J�ȳ���!��K���ۗ�'��1M(u��D�3�6�[e��>�D[[���Ƴ���1�1��WQ��@ �u�¡H8��˩�Jȼ#	�C�sY��=����O�h�{1��H�p>��� �mC0�E(�3���e��bq�тr�ڶ]L�9��L���Ht�ڴ�2�2��\�Ⱥ*I�*���1  r|�����7~��!��)I����wrp��Wz����m
m�8�Y�x���A>�:�KΝ �}1�d�J�K�	h�M�}���
�}�8�;���9����Y���F��~v���+ݠm:|�ٳ@L����&�M9�/���<��tT$�"IN). ��_a��\�g�{(�-���?ñ2[�HDW�O�����J��5<�%�\�Ю!g�j��P2��8udշ�L{]y��\\r�ǳ��ƥ�G����ui�+������F��?|*�bN��ŝ�/���gm��!*S$��U��@f��#���O]P���)j�i�A�d�@<��Y9����>\�َ̹Xfp�xT^��)�B��V׀h�.�g������w "\<���C��>�]ՙ���?l1����Bkki�t$KL��8�LN�5�k��Ԕ�ƙ���d�\|��W�˪���]Lu�K�����2����H��w6'�Ol]����[0�B�|���Ε���ۘ���ЪA٪���ēL�p����s���"��T�n�FC��2�ã����zôO)b����s�]u�ʎ��Z3�>_-�s�����w�˳�3=�w�;��f3>�X 5a�p,6� [Oms����"�疀]ұ��@,6�_��AJ�t]�N�Z#��@('��A�i�ɾ�ɹQ�C�'�m�������w�.���%��>��W�ƃ����������`��m}�$�v�{���lY����}�����w�I���e\<�1���r�_�E]�p<6�ޡ��wK�
A?a�}�9�)Y�횑sض�0��(�m�t�4P"�3���)��|1�K�zdV�p*�u���==���7�GI�@�������a~�]�D�O�^�+����CsQe�������F��j���c�7a �7L�!d���NRn�7q��y�S��W���(Cl�A�e�r�Ś\ȃ��ʾ[�l������1��x�f�&MS�C�Ɛ$�__X�j2��O/W������Tq&�ߐ�����xj2�����T�L�R�5D�ֱVǯ	�e�