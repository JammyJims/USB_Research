XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����S�����j}��y�)���B��oX.:�U)Y>��f��G�sF��Wn )��oP^��H�j	�&Q�q��/�X8�{�)�[˰FVUF��s��j?�HbjO����i����
�:�$�ӭ��6���;�l��6�^����Y�E��^�sp����K�fe��
�.1X<�"�&ͽ+E�n����)0�����+)�r�8J�{���Z�R�;��m���+w�n50��sS�3?;����Ʊ���h� �gϭ(9��Ӈ�����u�zD^�
X"�E����z��W���]�G�m�t`\��8�j�����4f�oN���:��� .�T0hD��S�6��W��{(��-%6L��}O���?�DJr����/%Zx	c��bÜڈq���~'�Į�p�~�]:A��r,R
1�w`�!���:�����j�>gV�mH���^����>�W��;w�-�NDX�D)�+�R#�Ļ�C%M�a��K�^)�2!�2y,'ZӘN��W���Ǘ\I[�m�^��)%E"�7�L���(�]���/��<�	�x}�br'��G��c);��n��b�r[.�n�HT(a�1�r�/��o�c�X1����^��~Jfs��i��'���ڸ��Ν���U1�@�m�V�J"����'	������`m5#�R�Fq3W��#&Y!wv����X��^'�7����n��ǔle?v��Іk�*��  �.yu6�zE�XlxVHYEB    17ee     730��U������4h�b'W����X�Jr\f��]�Ӗ��l�͝g�w�7l\=ڶx��%���2���V�l�5"�IOM1Hw��m��d��k�r�7�
u��t� �|�P�Vc��D���b����V$��IM������7b(򓰳��jY��!���4m	�|��l��3�����@VwEw��"���(<6���:5�>;�K"�$�#rnm�U�NԼ��q0�Ӝ��%s��|2����:��?O /v3=�؄�.�,f	���/cL�"�8��uO��ĝ�;��j��U�E&Aq�q�>���sR㕶 �u��ڮևY�B)����Uz������e,;UgxN���W{+f��Ok�K��o|Z����D�����BQ��u� ��sM���7��|�`� 0���7�QI*?8�8:�`+��-��lӨ5^�vW�s��l�V��iJ�=ո��Ϳj��i�fh���~����TX�4��6QԱ��qc�ۤL�(���1?i
��z8�r����G)*1��yJ��mۢ�{~��])��3��e~�_I9P��{<{�?��f�z���K���L��B��<��35��{#n���ʠ�k�
�tB���i�9NH��sA*��L7��23�����I�jbW�B�\����N�*;��)d�k�u�����yG�'ΰ�j�'�����������ӕ�d}&/'a$\�7>�Q�N�q�w�.��ͳ��v|ϚX��2�N.�Sދ/��f�m���?f���g��G�L���˸�@'؝��9��h%�G�Y�m��p-�e`FA�� �fqo&|Їg<�SE��oz�� ��!Ta�^�1g�����b��/���:�_x�d̩����C���;����`�̖�W+����<O%����J�>,K�VIR���"
���QC�뙖E�xW�-R��w������4�q욓=ւ�r�8��v�B�A��լ�˛��|	���� r{��	^��[H���?)U3�W�p֧�B)8q/�_�� M'�]�ɚ�?��/��Lɫ� ��� /!d��(��Lz��W�	yi�ߨV5[����;�� ײ>[A�)( 9��6$�⢑��r��ף���ȏOuhY=�����AN;��%r���N�2
Al����vJ���}(�e�^>�8ͻ���X�u�&��8���m�f�P̩�vT�l~QH+�Eڇ6�'�I��L�+�(�LF�r�����֞ }��C���J�`�w��$/����0?�i��Z��<h�0n�Q@KR�L�&©�?����I�BDFi!���"}�'&��v߁�YH@Gh�~�a߼�y�%F2���_\y�dY�i����`ݼ
^v��T����۩::�%r�ObF��T��݊#BI]���&�7��K����p�Ø����<6��F&�g�� ����g� �of��.�٪2s[��IV42_2�)�ݔú����D��d�=�:|�_��i���n\�=�����,NT���D��+S��d��=� y�<OjV���G3���B�΁�s:�E�ZdA�z�  �	��+��e�%��
�ch+9ι��:{�OU_�O�\wm�]>ߠG�R֜�f�];ڂ��1�b��������U\;S��@cH3��%��v��` ��-P�|�-ʾ/G�&:�R�9��=�ptȌ}�EK��ea�RtR�tDí�~�]��O,N9���k�7x��6_���.�6�k�kA���J�E�Ӫ��cR���J!_���VJ�9��x�2'�:�����yV{�j����8]��B@3�)����p��+%�r