XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@m���;���b��ֲ��ٟ�O���f�j��rn���&@5s���Zr�խ-s]v=�W���^/dkr@���(}�T�k���}�����*�P�H!�Q�{���O���#g���n���	��7;���Sغy��Y�T�j��h�� k�3.k���IO��z�V��5�H�>��)��r�r����A�EnEN�x��	Jd&��|.hl��gjy�.㙭�]�d�lߺ�7l�\�`�RU�� �u%�&����H�f_f�rp��dh���&�Գ�j^��O4�֗�Y�(��I�f!������V��.�qukAE[c�:y�i�k����������hMc.-��)�R5����3I��F�!����H��-����GW!��f�cXFը���l��Dc{��ʳ�.��5X������t8Й����&�o����N��$���\���w!�8��
�g! �����TA�]�	�'#��-H�&q��A�Ι��PY�4ؠD$<䇒N�������R,����ـݎ�D3��{BC� =% [S����r50�����}Ђ
1� P�pЉ�F"O��@ 	�:!}��x��<i���E�:n(w���8������� �*,�$���d��%<>­���} ����ɺ��Pb����[���� H�/���D�J���D��M���@:��/X�G"��w�b��O����X'�ERM��Ibɢ󝅸O2܊
��}�ԏi!�hs|ͽ�f���e�ѶuXlxVHYEB    29aa     980��b8!�93��]�Hw҄P"� �37�����>��K���*?&�f �mb�,\7M�N�Bvǋ>]P5M���0�TJa���#�]�BW����8�'�- Chl�0]A
�}U�Ϥ5��s������l5�J��"�vN� �+��v}^��hO�Q�����Ψ�u{P�wh��PeQ��$,{����b�z	F0�b�ŊX=ɲ�*2_>3�G�	�dӳ��( �V�H�zްA~���`��.J���<�P��d��g��6�gކ���;��|�R%a���⢇���O_��m�)��_������	�
�5AP��I~N�č�h}��q���{�h�ǵiΊ6�mk��.�Ey���p��>"T%Px�S!E\r���W�H%:
���U*�(B��q��b����z͌� yr��:]�&�,S>[�����=���H�0M6v�沒��8�)(7�^��)��U�W�n Pc�`�;�<��I5P��f��:e��� ��y2~C0r|���6Τ�~ʷ�SF��X��h�`���r�f�j�@ld��E?3ŭ��7h�n-�ք�It�Z�=�pj��l|+ �����������}5H&PT�]�H����;,���脼�?�AY#���@�	(��^�sä
փ�*(�� u���	���Lg�.�u����h?>����E�<�]����>����q�&�u�l��o(�2�����w�6*�����rZ>u2��wөR����,�z{������U�ŷ=;k�!�h�b��i!}����y\[�V��)���"�4�8�i" �mx�~'��4���w��'��,6��˴r�=*7���Q�c�DfgI��)F)f:,��"���c��(y�`�%=ЪC,��k����#��̫��B�=�dt�����&�2ѝ�m��˵����LDp��T�on`w%��>��{r��/"+��KE����`>���l� AxX�Jsu�=?�G5�q�D)��qE�-����"�j/�^�������
|^�gOhh��
^I�˪jgT�_���`E?��h pW�qg\/�E V�8�Ѫ�R�F!9��lA8p�lJq$�{������Y��j���İr�r)^��n*2+�Cb�D��P|d�`���4U}�nrp�_eW�u��/�`������q���O7{�멸��$s�).��\�p�� 2	Y���L�~8��O"���tM �Zř/?�T-�$����xf��*���B,���9�P�;��&���O��Ii��m%(OѠף�����l�n�VARL3H�³.|Ԓ���+���՘��i:&�:=�Lp��%�,;�>_��Z��}�$�c�'��s'���Th��lU;��n����e������b�%���Y�ĥ���Q�����y8x�c��¨�'�g�u%�Z�.��UƼ��dJF}��Ҕ�J�g���LD�L���|�аrY�{w�+[=S�3���ͨ��a�)(�R6rE9o���x�k��(�1�o����V��&8�u�&� ����n�U�$���p��7������}�Z�� ݊$clL:D�ی#<!=����'�,|�<�q%��i����\��t��)�U�R�-�D��ַz1����3y��J2ۢM�1��֤ޭ��/��Ť���a��J�'TP�o&�w�~��rv�H4	��W<}��&����t�FǑC[�ڐ��+��E9م��Kh�����e3�B�__F�z�߫�"�#�h�'n׈���BY�r�>y�q�ӛޚ}��~�q�O:�],����h��٢�\P/�3X[5r�~� v�g]H�(�"ݴ���)��z5�-�0��ly�ጚ�Lxa�������)�0��"4JV�z<�VR ]���{(\�� �t� .:�S8A䟢��
U+2֗(b���jر��N��|��SE�G�F|08�ˤfy�)�R���
�p��������W+O3 �RW�b�d���o>�C��/��z>��[_U��(��|%U������|�̚�0����� ��cg]�mI�hR.w
D�����߅X�7�?�JZ��s��j�XѠ�٩nn�ȯs��^�0X��-}��dZҢ�~\�q�M\Ě���@c�րG�7=�jq��o����)��{��L�x9,n�r�HGI�Xz��z��x��^6	�����{��{�1��?�>�U�"my;���kX1)ms�f�x����Q1U*P��{_����E�g��lѥ�7SS��\X�S |M���YxΗ�-�����e3���u��s�HI�"���Y^i\p|���-0�Y��vᩬ��gζ�vsR^w���m@��H��5�&&�`V���E