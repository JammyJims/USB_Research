XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��TM�����>Aƕ�⨆��ٻ��vT�g6h}
�:0 {��!``����V��"V<�n��y?�_�-)8�N�_^�m.Ę�5cVOc��B���h�ߙz�K7Ԛq����+lg+u�OܧZ�R�yP�;�\��G���@�1_fU�����߿��,�����%X��e�Ԟp�[�G��(Ɉ4�W�}�ER+g���v�  $c�U��`���8(R���9�;{��0<��+���6��W\�^�mpǼ�%3Vc#@F��?�o���z鍞�6O���\�D�V2 ��Ùm喔ɳRNJ	�e�f���B���Ν����T5-(�!&}�E@��@t���+�'��t�H���x"�v���=�rx�yI6����;���0���)py��~����`v_�qy��碨$�'�/m����OA�F��B�3@uzezA>�+o|Y��N��I���un�;l�����P6��y��J0(��mAZU�-��ֻ��*�I�
5q/��α���Z�l�\cT��_�IXTa:� �J@��_�����aJ�[��R��`4�����(��)��f;"�H0��٥E���^���A��,��X�E�$��kkW0H����K0A�(�Ú�ΑE_����兇c�����}>|G�/�/6x���-)�KSV���Du�1]P��� ����	�I۞�?W�E?��g�9(8�#g�kc�\���6�@2��*��`k�e{$gF�w���*F�MA�� �=����Y�s{�iXlxVHYEB    4885    1380>K���f.0�pPu�"��v��14�KdJ�07���q�X ���c�3�����)��gڞ �+z�$�%,���ޙ�����褅c �V�X�syu�y/�o���ǳ�$ȕ�|�C �3�{���! �pDd�����Yt�k�-�u܁���,\:�|�KG� ��r%�p��m%��r��;�]�g4�'���0^�ߔ�c�U�G,!b�]��1׉�2���\`�F�h�vX�Q���	h�e2�}�����u\z���dbg)J۳�K\o���~[�i�W����Ȋ�qż`"�>�cQ`���ꮃr�5��~lO[)��gЯ�@���w��o Q8�"��"�f�� ��s�v�_���;kb�ߑ���uh�B;��	?��EB���_�N^�w���E.��qfj{f�*ǟ[�O�p��!N�pnW~�r�\��
� y�a����>B7������8�r�sR�B
cɭ���U�����AK�=%*�6O��E�>��~�:F��q|\[�T�~�s��g���Ly��!*�S�	"���sP���-����P7��m>ie�X�HXߨ����6G��@&,�߯���WkV�o(��_k��\v]��*�=7t���.I�Y�W!�c������0u���anb�|�q�7ф��H�6�tI]�9R>s��-q0��S������C�[�98J�Gw�F�,�/؄u0`��@�F*a|�'m�A?���rt� �;H��z?�.:\$v�d����H��o���m���o˥:xoy��e�a�K+	��\�ߒ(UI���i��n70���U�p)~B���O�p�ǹ����6��`�`bk����Tv>µ� R��n���4��xZ�
#��c7b���ݻ��EN��s�M����DyF�IP�jK���|Z=4U]
JH)���g���FG]��܇�T��h�(���y�4=p�L��o#]�����|x�nNqP�с����p��+��];<*�w����xP5�whc���K!����=+��Z�0J��o�yl�Z22����ץ]i'���Du��G{fE��a���I�/ʋ��Aq��d���N��0y&#�
�fU��m\Rج�޸߶B�����Z<�!ݔ����u&��~7{f]�h�G#��/��vUB�ç���<7�[�BBN�p�H�`���w�8,�yP��lJr\��v���Nx~���E�ˣ�i'd�U��W�� kՍe���g�wZ�aJ|�v�zP2C`�	�Ļ��MϱSo̗��ro�v�K�=d��#�v�cП�&�|�+0���@9$R~��*($����=1O��`8����s
�L�G!P���=atN���R���K��O�҇P`1X{��p�+�y�'o�h����q����q�qXX���$<T�!�ݤz0+�|���ǅ�զ�͟��ZnFm�QĽ%k����ݣb���]S��iK����J4��xJ�7G�*T�V��@�����*fRS��������G��5W=��K��|v�'���G�����x�M��V�/;hA���|	&7b>ޘ�����4>�$���
g\�����pMܲ�{* /��$��dZ�S/�YY=��'��x(4�Rw`���i��Z��S�IN�$�A�/C��Ȏ<6�\��ʟlr���i�ĘhN����a#Y���ю?����G���׈wmq��Ꟍ[P�� RW�5�?���f�E��^�p��<(�^�]>��i���'-�3�F����|�7���ia�*X�v��a	��$�iXo4�݅oA@�wT�L-��b��d��pN��0a|H�z'�u'%̓R��z����x�<�;m�K�<��o���zHTA��2�Di���>�t�����Rx��	�!����'"Fx��c}��M� �$>�u�e�N^7e���[ʡ��x��)�>4d���D����$B&���"S{�ش�����n�pd�f��J�;;�� �3��9����Y 3����B�6�Ƈ�E��1��!���!"R��4˃��:���v�6�g�Ui�\�3f�O�O�@��|ۍĮ�|�k�E��Y=����Io��l��t0\
l5y�V�h��E����yz8�]f[oV5 L5�Q;���a���x��<Ϥ[i���lǥz� ~�pn���t2B�0���=��K��5(�����ܫª�~?짵b� ���nw�a�h]������vP������!NFG��@F�%���	��f���bi�ܛ��X��}o�K8MkG8��wV������]�uӥ�,�����1�+�r��n���W�Z�2�r�a&��������4|h�Ce`�,'��l�%%���"�����
�*����f���A�4�n�=7�u,rN��J�gRxT��+Z�@���iq�5�bi�V~I=�4�?0-0�s$-�˹� i*�.�2��qV��L���b���q+�v��OG�\��� �CՄ�9�ʨ���:�c}֦1� W�[:�?62W��9o����X�sC��']�����m��8���1��o�}�;7[�h�E/��*yr�Yq���v�iǯ�5��Ц�lڒ\���4��)�;R/��:F!��졠��Zvm���VV��_~����rArf�0�߃�a�D=��^��{�M����F�x`&]�#�|��V+&�L
�w}0B��v�L�����m�$vK�df����QъL0��b��E<>��z4�m�;X�J��g��[�m��4n���
l�*>�����G�T������uDP���d����0�r�$T��k&[L�Ë�|�
��m}b��� U)~�Pp�8\$�X審���R]f�ѧw`E���*6=W�~�ծ�'�@��������X2�r2�wG`�p��x��\�.׆$�$�qy"ɰ?/���==���}�ǉ��v�w�%�d���x��c��9i~J�G��g�]�0��jk�D��n�������?������܄��H ��I}w���Vp9���_�pz�9�ş}c��OAm��X��b���qi���z|�m!��@��źu�Uzf9���	�_즯oz�oV�F4�@9�2��R�Y�Q}e�u��Ӿ8ׁ�Ϯ�Q�t�J�X`�3c[5��������X��Ϝf�9���zd@�j��{D9�n�+�g��R�3	����(@��>��Q��1�o�xq߅z^�"�Q|�4���Y�{�h����kJ��$�t�n�W�YC\N9�$����SB��J��4'fF�zU��z�A� 8`!Gu܉���]��P����e���;UO}%��\�P����MY�ز�ˉ#�cD%`Q-1�'jl������x�;yl��ّu����_�"C����/V�0��xǞ*ŐB�˟
<�j�BI^N��<��rгP�}y�#�[r�Z���I�Tz�ZZ���s`�sK#���`��q����S˭������c�ҫ��N�%W��c�p�X�2��������r�
�����S��=Y����u'@S ���3�6I�<Q*#�e��AA+f�u�Y���ZJ���g�o&�8_v-�������*�~���[6�]��A}�1�;x�	��"��J��L8j�^/w���H��m&N�R���-d��B�o��{n�~���|�W�q���_J-N�z[��P�K�!��:�����G�Rb�N'�I�f)���,����E�:&�Ele�[�Լ�Υ�hǅc]�X'���*TTP��[�-7�^�8�NP�T���Nޥ5Q�Ô-�&�0��z�˝܈?P���ֿ��N4�2���j����L-�Y��4c��.@ň#�g�xm"q=h�&v�5@�e[t1uQ4���FQ�JM�}Ђ_�����d�iv�Ն���1dR�#&B���Bq��g3(��]�b�|�+�ڦ6։������L�^4%��!�a�rv>.��1~�3�3ۣ#G-��+��2���g�1� (Xd�Z�T�czA�鞯M��Ɠp�I]�� ����6��m�G�d��T�:�Ɍ�6q��C7��0��EUټ���X�	Vg#T:�fԭ����Ia�����x��p��*�Z���ͩ���f�f.T�F{��sE�FF��r�(�[ǿ%�� �7���N���3��2���Ŵ;�g��V8��h/�~>�niD�P�s�b�Ԙ�Г�s4���Q�-a����d2u�5
�}W*o2��^V�BN�:����(�Ve�iY��*�[��(zg�&����<���� ����>�L|����Z&�v��=��%���"R6M/#�#f�`��0�u6ez��O=���">H�ye�izW��Jչdo��4dh�h�K�4�w�=,T�$�)!�YIq�ex��wpЉ���&XՆ��?V�0o���f�k)��!�ڈ,`~��&XR��D$I����E�%�<�K�@����:�K�v����.��9�!B}��f�0g�w�g� P+ׅ��	\"`` �l=*�����K����Q"�gP>glNkXKY0W|V3���h�Og����5B��>'G��4I�t#;�|���{��(���ĕ�r������{?�#^4��r5z!�5����Čˊ�/_�)R���h����~N�x��]���Pq/�X�ĉ��G/O0Fr8v�V�0�������R/�S|��<����p��{T?*�J�'v��dE��[�������ծi*sd����z�1�^\����֛�;���^.��V-�,�F��xfc�R?�d��5J�G+��ɲ����v�5n�����Z��ً�GA��{o���㥯ZDw�(�dhC�yOӚ�7U#Ar���.O!��:�°8}b�*��i >=.V ����C��6��;(r�z2k&*��~#�q(��glh����$�