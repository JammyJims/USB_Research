XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����S���RcS�b�*'�t�(>|�ASV�)WSt�`���:��kr'��gҺ �<)k����O3�\bӊd
v|���.6���16�kL^YʱwQ'|��򀴬w^�e�-^(��	�	���=;�w��� 4�ʻo�S����J����9yV�Ö�Q�3`;�0�p�V)Dg*��ޏ_I���z0 ���NU4������pO��5"�Kl�)�����wnsX��	;d��Oל�.+�p�l'*�nv�LZ)`b�6{ql��d�[i�1Q��=}2v����9:h���L�O�*�o4�eҞ�pz���CӤ (�c1fF{c��O�EH���y���Y�gBf��%��ヘ�*��X�Kn����liu�[����� ���6:�q2�B��'m%i�У�A~|��N���:��_S�n�,�}�q��?����{��-Cp���1Iy���T,��~ ��q�C���5S��ă.�@�MB�R�G�MDe�.T������F�@\y����p<]e���)Zxɿ�9��$"�^z,��|A~�_9��P=���3�����xT�y$�?1��w�Pɒ����Hf��2{M�-�M�<�V#(f̴Th�{=:��7˔�?%l�'�j��gj��gZ�QNY���LX��c�f!��!�P�����{�A-�s�̉
����)�=4I��aUYǂ�Og�k�x��wO�B��~�%/
u���y�I��R�J��[A����৲�>�+�TXlxVHYEB    4459    14808練���rG���~w+us��Ǒ��r/[c>�W��9���Dгix�
1 ��C��Mv��C�X�ħ�5�� �܊X6Ą��`�3��^�=�)r�?���_�I7Zט���)vF�B���ߎ��)z@ZoMC,�;���^�gGm�^~���u�'\�A j�gc9���ut��o���+���IT�kJ,�S�B�G��c ����tHBt�nVC��m߭RnL�ZkN�r�
�e֝�ܔ����1�,�זDK��h$��Fe��7�+��0�d~��r���
������M���[O�I���U���?	~�f��L�X�Qڋ�K���{�	Q���_(,ዣ�S��NC�}����瘞��4(�z�cw�7b5�RO�T��S�o�3���>������'f@�߱e����(�1��)ד���$��t��<���K޾��ɥ7cJͻ�e��GW"�{�YqI8��o���L�s�� uޔ �M���H9�8lI�cr�0����v��d#/�x�n�­nz�z;��U]�@�7�Xҫ�)��Wc6Q{�q�%H5:�����b�{�ls}oV�P��p�mH�d5M���tU���?b�.��Ǖ�����.��dk�<��{�qQQ�"�CN$�)���~\��u^��{E�m{�	��Nt�Ņ7� �~�l�QUX�mr��*9�"b�ٹ��H�:���<yP[�lT�c��I�&*�/Iov��Ǳ� ����؅��KXF�H�]��x�/�}[���w�kI�kK�\}�#�MZU^ڶ�"� �`�myN���-�ֈ\�:�=fY@}��s@��ӞV�lr�� 8��8�(S¡8�Y~�oOA��*P^�e.��}����f�Z���i���@iFG��R�v?�u��8�u;���#�����SVN��'A�����;�d���?�0���\���W~iq���4��އpTB����m�g3D�~K�])$P��ŗ�+�&ȫVV]-�BT���������W��J�'��?^�E���=���S���P�������w�
����ϼF8�E�K���Cp:�ڀt;a��Cf�u�r0Y��.�Ve�����8jgj�ɲFhſ}fN�;��}�yL�L�1i"��ЊS�=������s�E��6�D��X�ʭq ��h����+ �[HTV�ۆ����e>��j�h�P���j�J��6e��1���]DƩVL���$zުJ���|�d!t�����Ȕ ��h����\����G�H��f�S�z�
lu'�ɪ��L���K#Ӟ�/A�X!,�Rks��M۰P���̞�y��"HZD��;�r��+!��Էtv�=Y�#+�+U�ǫ��?{��Ē?8U5���e���$~T>`�<�lRv�jD�#�]�Ѽ0z�R7i�*e��ϼ��B�|��g��"p횚���(�V(*<̿��Q�1Z
�u���1�L�e������JS3��I��}�n���!�@�ɛ\�̵2T�o�_�k�¼-p3����>�_�0�U���-���,��j��漄>�mK�&#O����R��~"}�]aVmٴ��Yt��B4���n��|��PT�+����{�Ǵِ򔨉[����1�X�HaHwcy)U>5i�LZsXItL���V��GgF��S�-��S�0�U�"��c`'�#��>����Ɍo�j�]�86�~�Gj���^�� _�J�$�~C`�	s)��+p��x����n���}ZE(]��L�&�ggW$Ϻ�~����kE�[v�J��l����l�L�����bm���gj�*ДHe�d��U�S���?Q���z�ȢO�Z�n,S�Bƥ��z�s.�o+�m��i|�;s�eij�/)?B'z�z���04�:�,g~���� �t������W�[�
Y(ɕ���9cz�p�rJ̞�$��N�� OY�c�#���N"�:��t�s���r���:(k4�Dz���݊y_kF[�4k�����i�$�{�>:w I�%���)9F�+
����R�'�ҺNԌ�%�	"jD��bڬ\���sH��)�	��܂P4S�r��?|�`!?;�`�:�o��O�SW�2O2U����O�r�M"����E^�qd��:r�)��ۧn���<���Ӭs�_�s=�j<7QFs��1,i�j�*Q�z�\v@�K=!�~������Ô���w�%8�*���3\�q���Az�s��`O<��XN8����J��d�TS����\<*�j�(�Oz��䬝�4��Zb!����1�LOB2����U�`����c��D?�W��~��Xs�x����4�pe�3�C0��0��c�>��(�b��R�`e���K���f�2kR���S=e�ŷ�4�|c����W�Bh�!�(xJ�%�:!͕�Z��W/(���Q�[��ڃYb���@��1���4�M!�"܁��g��<�V ��nF���L��e�Ұ�������IkB�r��呞tt1J��V�{�b��]:-��ˡ]�H�
WW��J����ȵ���}���s�T�X9]���*h	qB��րA
����bu�,���E��	���}Θp)p�z���U�1��'�k�Y��g�솃e�5.�[�:� "�_4�����1�ba������ZE �\��w\K&��k��6���Ŧ_`�5��2?��jd��U=:Uk��x�HeR�r��~�=��T�2̊@X,�~O[��%f�j&V��E��>8�ZXc�P[~�]�t$Ԛ�������y쎜;���[|�3��<�@g�u��*;���U�����y}6ZuCP���f� )c����������,�I̊<�.��$��tD.�Sqd�T����~&۶`�@M���0�!��lZ���h研���.Q�F��d9���O�F+?<| �цJG4O?k9�Iƥ���\�u63K�x�t7!��Ͼ��Fe�S�n�'��q����i��&�� k\�%`m�fI�rH�����q�� 7�p��z�Gk?��m�G��ȵ��Lo#la�1יD5�cx�~
?�n����`��M�6����Ծ�_S��J�t<����Ͳ��#����F-BE��BI�!*
!��X���%�#�2��3�[�k�4��:��?f�^xօAI��Jv�z�D�l�s�[�9�?��Oy�7���8U�X�-�&��^I�M�˿��� ��D~+Ry- b
7���,wr	{�~B	�����mKҗ�
�憛6�o�錅�{���Ҵ%��[h��W��9�$̑:u^h�>�:��·�-.y� �)����E<���^Ȥ�O���`��+�<{*	�7�����7W*�7k�3w̛�#D�mX���{[�?hr�c�談����'/�Y�M7Cpd��ۓ��cZ��$������f���ʳ��'����������L@��h�772���؆������U�:��-3�"I) D�>��_{Y!��������q�\t����)�1���Q2]�w@����4������^T��s�>��ђ�x�՗6p�A5����͛}�è����<��aL̈*��}#�a�A��m G��9�l�#?ۣI�#��h�=���7�[ӝUX`0�\���2���o��)p��?�?��A�D�ҳ�fD�u���ʩ<��n�T��G�/�3��򠻽�{n"��d�4�u��#ܕ�@����t�:b�h&g]
x����=�(�YZU��:�#�|~-v����A8X�}`.���j��|k����\d%yZ�V�Z�
t�\��Ё�J6�f.�VEs��3�9߂��ؾ�dc���6o!\g�%�)�+J�m������D-�8���X����4��X�b�SƧ��F��v���K1�ʥ��f����9.~!v��jz5�*AT%������!Y����q8�������:_;�R���mZ�h3r����p��֤g�W!*7jl����f�a��!Z����y8PL�.~��1�ˎ��[�H	cV�ډ<�&!���:*��ɜ���sa)Z�pq1��
#i���b>1�d��gf66;Gڡכ6Ѐ*��8<+C��0r�1o3�J� Un���:�\��~�Pێ�
��v��2���!v�n�xi�u�3� �\1w�#��(���мP�����bꦻx�&�1�2�5B��q����I�+
�p�O��_�Lc�6�#~{V?�����Æ��8���2�`�9�G���c�fH������K�i��`4:�8ڥ������N����8M�_���eψ��A����@�T�j#�'�߷"%cJ�&�Dm�U��������rsi�HXpk^4CL�H%4��uQ�Tt�:Q��D��/aqއJ�6���
�eF�N5�挕x�a�=��e5eo�MW*Bo�����P��'��w8�[w�N6$mkX5� �2E�^~��	~6Sqr�o-n�[�����Z"%&^m�{��w	f��O����nR"�$F�����ҖIAb�?�z��*�k;��9��W5�X��uN��� ��$_A����1�_���J�I��Oe%4�/�=��Y ��]��G��f9���)�G�
;�d��0ٗ#�L�����e2��xy[��l��~7���B����eS��w&����Ȱ,q0���>�������W&���^pQ���K7��A\>�S��djwt@���!�.e=�2�M��`l���z��0Y� ���d0�h#�CN
g�ˠ-�1�t�9J�	S�U󤇋��~�=A	a�P�̝� y�A1���|;j�$�D>S�H�Z��ޡ�g���E��<j[�#;�z���'=�,��5��~����V�F�x���q�<�lE��F���q��!��#�T��a��&Ь�=T�RL��r��`�i	�j��4���}߈�گ$+ �b�Y�e�� 3g4K� �o���!V�ʥ��G@�Bn2�3b}��98��*�	h`�эeg���?���Gt��ЎD��߸�߮�Ȫ�\����d0Z���gQ�v�c�����#l�qLwY���d]#����7:�Y�^���l�����c�^�M�Kn�k��d�&�sgx�,H��r��5Hƫ���h��uc�+�Q5���"������F6M���@"��r0��%