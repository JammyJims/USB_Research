XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ב� �j-�/5�rS�w󠚁GH�*�?u\����6S۰A�% ���0&��vs̶I�'7�|���;�QQ���[�a�7�	��*�?b�L�X�#�]�T$A7 ����8Vx~�ƽޡ3딠�a}�d�4)kY(��ͱo�����yDL��S:EBD8�0�`�;�Q��v��eF��\ֆ�_��څ��G$ ��?$_��u�F8\�3�[9N[f�����܀��M8�Ş���V�n j���<���K��X'�3�v��j���E�:B��t��<�y+-�2��4�.�m+N!]so�zU�J�>ŝ8s��1P�Cdwߌ��Mg�rZ�?l3<~!J}��� :Cn���D=DM4�`{u|	_;�{��<Ǐ�h�����/M1�;��P�T+t{��|�g� ��s� $)"⟂i7��(u���ĵ��C�]�h��+G�v��9"��)M�yN�ٗükwzUn�Ѡ����sV� ��r���Ҭ)(�\W2 ��qށQx�K��.�yg���:�p��5c<�[?!+I�9U�-B?���HS��0]�"_5Z��*Ƀ�E!�V��Z�r�����M�"���0�F|�Y�	��g�)�@�j�
�qOw����i�/8�C+�JI��-4�&��ʺ��)�܀����%�gw���,�q�tB,�������S��nh��-3\!�"�c��������-�����Ӽ��2T�9�(*�&�X������ ���U)��<�i�k*�UXlxVHYEB    ec6b    1e10t�Y���"v~Eo���+T^������|��Xt��t�?7���~ֶ +5�Hip*����N/�4��=b)y����b��e�"[}�/�+�T���	���}��>��b>� 6����g��^��#.w3�M��p��ұ�y��2�j�����bE��#"�G�|� L�\[�I+�_��`З��{F[mI�1���0��H��,�;�<�t^1�Z�@FP8Z�0`"��К7ݗ�Ҵ ����,���bh�v��\�'�'�^s,F*����d5���ϐPYE/%���{��=jowHǸu�{�5r�8��Y�9����M0qge�Q���ߧ_���?7�0��! djDw����J�d*F"�(��!-�E{�1��h���T�x 9`��¨j&����w�2m��t;��&�PV�𢂆�B	����i��/�(�2o���Kyc4ɰ�n�'�����c��|�[}��^�>��rZ  }G����)��-~!�����0{��U�?^�Z�Z�7��VF��`����l�D
��{!~��y�%JO7M���yr����tFj�ь�������6\V�����4�\qڝf����n�e1���Jdor���?��,����51�D�O�E�]�O���/���6`��]R6�xL�fh+Q`��&�Å�>U���&�tO�H�ߠyIￕ��T��<]�8�ߠ��@:	ҝdd%�a�������3�Y>�3Ɗ��6���˓_����XУ��߉�27��}���Y�L�q����1?	HcY�G�3��	S�Y׸8%���tY&F����<θ�$�����]�?6�Ԅ���Wz�f���a�v�y��nQ�Z(;2�G�mO%/��d��v9��ta�]$�.�*ɪ�
fЖ/䚶�~߭�� ���&Of���Wx1�����fR|:aݕd�4��x��G�'A��,�,������{~5mZ�[&N���T��<'ĬL���#\(-g��Z��OU�%&��D;|����Dn!����5��G��(�����dtN�/,V��h^ݠ�!�������7��:"ϡ��DSX,���S75"j��R��>yͳ[Vq�;��	#O������eB�������Ӷ:�p�kv��P��#zEpϡ�TI��}38|�R(ՇN���JIxҫ{+I*����`f����<�\�1]���I��1JI�'�G�F�,%�OɄu@��/�A�uԑ`�$�������}ٟ�R�٪�2�=<eP�v5���E�\��㼂v��*R�J��s�����0� cㅯKGr�'��Ձ�MTV������;�����y�,�s�k�x��ɧ9��{�yC���I���������~2Pp����|���O���UG��:��ްDEv+��)g΍#��H����4�|9�y�1/ͽ�E��ө� �沂Xg��6`s$yY�+AE�Q��d����(��v�8?��w*�D��y�k~���Z,�c��lb�ay���s���PE���DW��~�����hSܖ�H�\� ����5�}�)��@!In�E�;�Y坕ښDZ�8��},����
Vr�Y���������uus��R�p"�&pc�����Mw,�<�6���٭����P}	�le�a�a�RL'ۗ��@C�RL�	�W�)
�(dA��č��՝N��5!Qs��r�k\���eo��m�t�F�HpE�,��p�a�8�U�[%�	o�'������*� z�/u����Y	�R'p��1uD��"��/v C�2��6ά&���FQ�<=�qo<���dy�2�0�^q��8B��Ś�T�ˍz��0ғ�c� ~�,O�)R�
�!<���t���6��+���A]f�[���̘<�(���i�
}A��# m��O>�9��$y ��2n����g}Fl=�3�U�E�Q/�I�WV g��q`�'<KR���L���e�	@㛹̷P���Q�ho�;��+�[â�Is�?�l�6J�{�������H�m����Y�8W:������/�6q|�G�U�����r��#ߡqB�,��I_��R��щ�[R[�������=���t���a�>��C�6�û*�z�(gU0I��w�k���#ź���py=�5t�W#���<�$�N��	Y�x��85�a4��;u��Ԗ̹��'B��o��zT6P��nn���L��T�|>B�gdN6'���3d����J+c�Ag�mQ��``�0���@Q�2=��a#�JJ�iD;2����F�m�Ӧپ�1 S�&�2T�(!�x�y��<��&@Տ�J�94�;N��]�)XcT��ՆzS&�ba>a�k��y��Lv#�	0��t���z�n��޸�a�Gdz���� !����i2l�`�(A�S�.q���IT&! �"�&Qԏ7&���:�Ѕ�aNCaЗSFW��t��)E!e��1t�0�ܠ_mb�1��\Ʌ�~�q��&�����CH���њ<.f�I�������?go}�T���k�^�`��.8q��;^fY�!�Iiu]y1��>�7b�>�j3!H6fzL�}�%㶯m19@���tn���C
�ޥ���I�2 ���T��D�O�3���)JР�y�'���g�DtqA���͂S����q����mT$l���=�d�$tH�7�S��GKe} �4Ū�@�AXcE5����Uc=�k���^ޗ	�c���.�s�.��C�(��8�D~�>�I۝�J����� #�F}����Z���-l�@d_��v�V���S�K�-�*�͡\���ɡ��B�CoAK�<+}#p�$��_�!�>l擮�@k��Z&�;�3$xhN�1���o(�Ծ���Ǟ�xOX���a��fU��z,d#�ͳ�Q^ɬ��7 �ۮ(������X���o�5xO�D�������g뮩gtEe�����IP�8��#�ז�;�sTc��NVC�e�]� �txf��m���A����]���7�F�9r":�W���e%<%9��z��}Éa����ղ�1��R�z�]��K�|�˲���>�X���H�x�� ��Uگ�gXT���_<���Z$j>��j57jD���{�u$���&J�d:Ƴ����]L�P���K�Qf�*�6��aV�hi�ݫn�$��eq�zMz����7���� Jt�H�޳��h|h)*��c9\��������?n\�����D@#�P@��-E��OP-�ګ(g�<6ʲU���޴�y�7��$����Z���w�M7y�mј�_���A�,m2��<X�b��*A���g_���aQ12��fk��a�H�W��b�d�I5y�ex��9mW���t�(�e��^�	��9���s�p�F��μ�#����u�7q���'Lf!2�6��ˍ�Ž�����;{��􋶿'��k��/���E�h�?*D��0��jYY߸��z��?��*�4X-���!����2{��t-t���_�aݠJ�A
�X�7.bP�PG6K�#b"��/�U��Ռ�\Ϡ	`�oL�g�t<�bm[�� }�˨�}��%�'��*�v�6�#Y�_�R�=�H���)��R���M����@��(�TJ7bF�?K�a��s���d�(�D�ֿJ����o���1�mN�ˁ� 4I�6�ncI���n�X����Aa��t���&ϙ[#�-�8b��k{M0K�:�>�!\�3�pu�ET.fؖ�)�/��� �=F�̿��
��T����k�'�H��-r�\_�*$'�K  nB�5�����^ۥϩ��4����<���y���@���Ub�&��>z#1i`xZ��RMx{.�B�d@>0㊶���p���j���>7F��NЏ-"���r_�����i�z2�W�I�,�}22J���%J壩��w5�;i�M�0�?^1̧�/��k��cXc]�CE:����$�ѝ�.:Z�3U���i�v�i��H1&~z�5��CFXW�3Uq1aVֻY��'5����5Tq��͜M¸�>	#豱#Ax �_���x���Z>����Wk�˂j��^��v(jҗ����.&�P�ab\;'?q�m��A��φTVQ20�j��=�I�S�S��Iw���nS:�mt�p"�4Ah��tî:p��y|�C_��4��z�6[I��	�&���3�|���\�l���T�2�g�7?�qQ�]�Z�qt+�q���w�^iC��@��O�TI�&���%��k����P5I��$�窺�q2^�D�u5ti�pL�/͔t����(�>e���6u-)5W�F���t��j.bƽ/�`�I��ԁ�:�T,�@ldo.c��)������v�D�y=��F΄F�~F5����>	j��nƺ�K:v�Zd絫�@���A��#;��F }��w�~a�^eP�Q�`�i*M�8Xjs$1����O�{��aΎ�
PD�*�ڬ�4�lC��v��RΙ7����atF���z9�ݔɘ4��������%�ic/���3;����_���2jX�qX�mV�9�P�����j�3Ι�Ŕ$n�	��.Uji �0
|ᑉ�=j9�eI���X~t��&N�?��t ��&���,�1�O�>W-��ԆR�=[�`X壹lQ_�@j��n>���x�Hd��<�Q�X,�)�k�R:���~Ȅ!�s/6a��˰�b�����9_�?�C�3����IH���KLE���@��'.{���}4��&���$9��d��hA�|yQ���%��1b,�/zUV%��.R�4��K��]}ͼ���@��\��0P��g�Goe��$�)�3�X/߯�o�8���-:v'�s��I�)$�IYDU�����	ؘ�	U7�g3/���/Tv%C�v��l���O��[[�X�����͢�%�9�\A>/��]@~����аM��9yу��K�f�H]ug�МlZ
%PUK�:�h�β��V+�B�"s*�:˗g�5��̱�V�Ȕ���2�̎|��W*�Pɧ<E��	ƨPГ������pN�`���!^�C���1w>{S�$�����[@�a5��^C�{m�W��ߨ��е*X_��I0�"���5XmH��>��1L����Oj/�wڇ�&&v-h],ũ�'�AF�O�͔�ȗ.ka�TDh켞A�XZe���oVP�3t�{���B`���?ͪ��x�tw��eu�:+EҀ����������|�^"�!k^2�h?��3�rꚬ��wQ0:�<��Z|�=��4T�"ۘ�M~Z���;����#�TxsUI�f����M�pFZ�Cq��8���H��wL��w�����!�զ�K�)0V��� ��8�/�:p�EU�e,|�Fݕ���s�˻��n�X�K�\���V�x���3��_z=���XjE(���.�HK�NRS9jjs�gŜL��&�y�!*��
�"3�YKUĳ���u+�a6(s}�x���n������ �0=�	0;�Y<�� �y-�4ֲ����ꎬ���q����,G�"J��,n�-��ţ��x�����ɉ]�,�DΖ�\��Z����}3} 9S��2�6��X�=-G�6��������"@o�ы�*Eh�W)��2�?�Վޣɂ�n�l�G�=�JXuC4��1�y�vH����o��e��\��JB#]��� Ҫ��5��92S\��24��Z
<�z�a'�����D{O_�;f��UWM�
I=��y8��:fh6����j{a��8(��#�_P�dsAXlO���f�� y���$�;jγi�	t����P�Qt��9Ô�f߅���Tq꺜�T��S�ݙmgu"�/���B�m��>~?�����¿��&���x7�]+�­�����j��:����C�	�
���j�Q��"T�\�7��X��Dz����U0��m�R���r�7��O�>ӡ��6�"0�]� �sM�X�We��X7!�����̘
u�ͳ����bHY����/���!z������R%%�sə�)��N�<��75�K�����DIjg��~�L��ҮO�4NZ=FfP�F�T�@_a��i?�g�I��m�_d|^�+��Q�������u�u��Vѵ���"(�"�D`%��
�ɪw�9��a!�>f�o�$�޲�ޮ���9pj���c��䉩�6���
<����_`xOb8��GTx9�*�+�������W��ՃȞ%U`TQD�W�L�v�g(��n�����TUO��<�qp�T����N��-XMʓޭ�c�%���ן�A7WWV2Oy����m�j]�hNf���5`BY> �@��Q��r?'{
D�X���y�bL,7b͞��l�1�Wpe��+�а$y��EB[w9�i��O<�P���(����j�<���������M�c!}�w>:A#���駭�
�%mo%������r����_>n<�E�\����[˚�p�N�)���󕾴eO��( �_@Mզ�b�uͲ8�B^��$�|���D"PQ�"4 I�v�n=����v�*�>�;4fS�˜neb�5m3)ҘT�CJY���e7�*|;Q]��Y4��Br�8'���i�����I["�E�?)�苦UpmV�`v�<�C��
>;� B�^oQK�����@�D+��r-�t~���ىBZ����k>`��}G�%s����xo�Fu�z��,p��+ǉ�*��咇���}YA�G� �OȖ�N�=$�<�Ԯqר�y�3�տ�k/��k�B�Z	��� �w�V���F�vg�prSe�����=������&�0OPa4������Y_���M�wǚ�B3f����;����C����G�9·׫�����a�u��ы:rN�X�-���<�_V�[o�CJsjގll9x5Я:�:��P�4��9��;����n��ϋ���e$@I �C}��׮�Ul�,3���Z�Ja���	L��s�Ӆa����G�����4�5��_����z�)�s���i�xU7��b�\�o���.㹩����c���(��G\�I�4���!(�U����y}l�����,�B��d*ᔬ�s}�X���ƈ���Dm��ʃ��7Fx-j����͜�c�L=�x�Z�c�h�R1>C`y���<7\.a��b��ј��5�_8�
��,���J�����F	+㰎��8߸=-rV9�sg�_z�zN���n��E$�`��F�.H"���ɺ�����Grq;s�P�*c��NG]2p�s=�IxÁw�>&#k���$��m������V�����\�*H�Z����
� D�p�T-xq�S.bx�;�r�<Z<�b8Ʃ�2?M�0�[�Ѥ괃�/"_`I�\s�c��X��$�$[J`��Ǉ�Ux��V[M�4-�#)�ekRwv��4a��@�$�G��;3,N�u7���=��Ε��ט���>�-�Xl���"�q�[�\Ov̝I�ѐ,̮����F��O�+�M����EN�y3��غY@�n�}�;�Eb�b��X(���C����7Cx�g(���--g��d�Yr�B�