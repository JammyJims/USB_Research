XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T,�0�Nt~̌�<@�6��X՜!���E���^���s���¯���B�$a�66^
�g�:�G	�5����>,�
!��zb�ؽ�A6N�M��7i:G�8Y2�� �L�2ZI.o]d%CS�Τ�jD�;la�����h1�x֑��Q*qy��m т})HK��9'�z��}%�4&Dś�� �����^D{F��2��xU��L9�-8&�o~��K���H�T.�m��Vͳq����di,Q�H"w���2z�.ڞ����}��Y�Kte�����H����9�� Siy�o�EUv��$�!�����n���_��`�2%�Jq� ��5��V��}9A+;C�f�i�5�m�^GF/�-�q�N�"m6y��n)\k:�r���~n������m�,���;�ۇ��qkD��{]L�G:�~:�J[^�'���-zZ����޺c#dy���r������	���9�X�������#�ד�ޕ�Q2��,�𣏋H��^�;��QW���js�|.��(�H,f��y:�g�y!�v.�"/-�K��#[�j��"���	����*uy�\� ���*+���{�{ O�������9v�������pH]o蒱"A��5~X�,:���mzkS;��W�>��L���_�D�=�K�8˧[��EPD��<�?�:����F)���A�J����}@�w}���(x=��݆����Ͱ����+��p;����YE\�,�^����ߗ[�?���~�U��
���XlxVHYEB     f07     6e0z�V����ܽ@�W ��:��}��|�Jf�'� ����&Eѣ2�:��C�y֯�]��ତ�fH�px�B���8@�M�$���?�2K���t;���<���2�@Ĥ(q���ᔛ�K��\��3�|VP��imA�L,�Z�p^&�]��~����(���狜z� Ⱦ���Nͩ��uۏIY~#�*Ig���E�e�u
U��r�e�t�zP:�\��~ĭBZ�*v ���J��I��3f��;rQ��,�8-w�4�3a��(E��P�p�u�M�z��f�P�q��z�UeA<�xB�,�G�p�g���鎖���_�:<>�b�	�M������x������)�F���z�پ��o\������W�n�1r�|�:�N	9P߾�b)|��Iб�}�	��Gg�������j�d�����b��F��'K6+�����F���]\Ny����1wA,�5O�%a
��i��]�7�sOv42Z����p��b��Qq�ER���ק��9b���:ч`�~b�.�-��+�)�K�*�O,"<L2����7������-f��nB�p��� h���}D��%�[`���%Sa���I����,�H;�Xh�<a�Ύ\���<˝��w:/��h�ې����KŖb�ˠ��6�(�Au�b�ˮ`�� o���w��(�j �&Oj�Pď�H/:9�zo��W��o�\#{�-�n�hYH��z�ۦ���_�b$����/	�� /�t�hݛh���_q� ���{�dp�NYA�Y2�l�M0G�b��N�Yi@q�5�O���@�/1AC�|�pk�ǐc�!ާ�Y��V>��n�ZsD�{-<����䨵� j�6��g�	��5)�℞o$���l���t|?��h���4V���v�R ��Ԇ)A�	�1�}T]y�)$Z��d�\�j8�`���2��rP-���]�r���`؄NJ�Aw��Y����������|�Q�dH�$�y;���a�V��E�{�=�3��L�U,���=�@ݜr���*����AgI�D�1{ ������)˛>���y�ۛ�������  +���'����'��KA�� ��*N5��Sbl�_����_(O�@���9�r�{PK^l�@G��y �\g��ȩ�빑�~[��F���� B���v_�NfV��~7��C���g`ib�C!�Y��A4�T���#
7�(�A�#��. y��)JŢ�I�R����v�}�>G�O�ӥ+��#�S��0�ų�|G��eP4O��k[:b{�����M���2�_��JQ�+��sa��=�j3�;∈�c��[~`��%`�����1}�\ÿ$H��^�D����-�ؤ���w��>7l���9�U�(=�fA!�U��K^2+�sf����lg�����ל�
M��_����7�;�c�Tt�U1$�� �шP��PZ��X`���B>i�$+��y�ԣ	XX��u�� &e-������{��C<�11�V���ÝeD��2�(j�>��z �p��=�g��U�-��p��w��ڤ�àO��/)m���fʓ��W�=��z$�bU����7-���F>:舡��T(���w{}L���<�J)�g��Ѵ�yU������r�V��jÂ����ꉨ���*.�X��z�B��	>sP��I3e&8@ӓ����Y������=�'2�痱b/��1i�