XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���F�x�!$�
J/F��:J�L��k){�ct>�bz�]�Μ�ZIZ���3��K̷ ��
�ߖ-M~:��0�J�U��mv�F9	��jvx��q�t��W�3>��cz�J�O����]������.W�@s~N���̓����U�Q�|C��&n�m��4_A$A�dP#:�}BzVl?�pZZ������M� -�-+���m�s�o����cmgQ��
�	1U��[��p���3���[��vn��_�gϱ�LQ�����5N%]��2G7:�����M���N?E2�U�s��4=3�D��Y�18J�ņ#�kB�ڋ��̨��=n�R���D2��뀵E_Q���2�wY8�/�H{�DM��2r댟k^�PP e���Y }�5��
7I��^�Jvy����bƸï��s�R ��f��`@��>��������Hâc�X��5m)�Q�^������z���7@j	�&��抜YyA�t�Qi��#]�r�ѿ�K��~�Jp���sR-���=� ږ��y��&��Ж���b�:��+xiş���ؠ+�e�����,�l�H"�z�r�g���j���X�O6(l��^Kx��[D���b�����˕C�<,�ll���G.s�S��������g��s=���eB��!&K��1����I�RA�>ب�?�tA1�'g<�s�c�ܥ?zf!@%y}ޡ�6�RԔ�F�����Z�|4���F�L��XlxVHYEB    2ec3     d50	9�Ӄ�� �,<c�d��S�ʒ:3.ԑ,��(%��I
�d�g�K&K��v��*o"I,����H�),e�3�u�1}�b���W�4�Bqk�9����e����sS��;&��0��[���g��v���|�}�{��Opc�͆)��O�E�wW	�B�Ί_�j( �@�bP����'<� f�k1� �s���X��;��5z��eA������O�M68��$�Iz�o��N4���C%�z����{�h��Ö;���#��-���t�J���q�IV��4�T�:�.2
}!f�W�
�R��Yۿ�9{���U]CݫZ�(g��v�(�c��;���Ě*���l�"��'��`�(��H��|:Ώ"n��XQL�K	�^珈���?�<)�5}K%5��o��
T8�E���Q�yyE��5�\�_Vqؓ�l� H�H�F2���:��/��(7��C��Sv��h*.Q;6ܝ�n�7Ogi�����!�S�q����'���y˰5F��nn1�����F4�͓�d����R����6ob�"%���|��?����3#�U����d:Qv��`��Jo�.+D��>4�֛ڝV^�����o�&~r}�}>�"x4v�m�x�Il��N�Qw��u)%p�O6w����MS�k��Oq�7n7�Z��,��>[(��5�.�:k�m�II]Q]��=uj~a(ɞ%N_�:�lI1�<!�b��7�9�օӘ%�:���E���f��Uw��&}��e�ǲ������m�M�-n��o/�a��(�`8%��hN�1�Mp�y�75fC�\oS�'W)��x�����(�uZ��y(11ᬠQ��;(f�a���N��P��^�c�Asx�xU��T�A��̫>s�!v+'R��+�Z7�ƿh�H�!��OD�#�n%���E��D�0rz�?�d=�	
s�Z���.���Y}�,�#U�Sn���G���0~4�E��22��kR�{����!�_=����a^ė���<ӳ�V�z��JM@X�b�e�}�%��@H6v
<mpԿ��f�C�	 ���^ɟ\m��D�_y)XL# }�H몣�����xZ�[9Me�6-������$6>�����p�����$�«�벌�f
�6���J���uTu���Ǭ����Ig�ٜ�Ah.�W��"	,A/}���̓mp���S.U�%�L��THm/��-k#��.������k}?0�������XytzV��e�Py~ch��^��	Ag���G�p�n[-���9�����]��=W��>е#ޞЊ�	�4����r=�G�"}�A���J�p��rH��~'��*�ů��M��]�,\z�'���`^4�d(8���7Ho�پ�������чnH"��d=�L�¤�ֈ���5�C�����,������w�"��fF�������ف��嵽q�:�:�q�m���֪��X�I/���kn�->bVN@���.0���s���r	C�m�G� �3t[���AF'��������|���%�����s�t!���:4���en��㽪 �W����K���x\�{=�}%,`	�u��a�p��6~l3E0���|���:g+�}��e^E�U_&�!чR��ǂ؃3��ڄ�d6�*������1$j~]	���Z�?Z�RG��ҍPg)/J
��E7�RB�T�O�͆�����;V�si<Z|o.Oe�Uϝ�zlf7Ϳ|$�S���[�	cWˈ��b��~/)��קCʖ5����Ԋ�Ϯ؍Sl���͊��Y�T�|�e8���A�����9>ܗ.�s�E������uY�7ގ@��t�{P�����t�3(2�,zKrY,��?I��f!"��yT0�^�N�/gc��̬���+����o�cAT��e���/��&�E�t�K �歀R|���[ւ@��c㋌�{��9TE+���X�`9FG�����ų�?(ڜ>�������1J�n��G��?(R�"����bQ8��x":�{�gd~�9@��h-o$�:^u� ��'��')E�%,9�=�o�/f���ǘZ�mhR]�dur}裞��&Ez�F���F���C����Y�w{��z�D�EL�k��p�{~|A�g�U��ve^�1/h>�ꔨ����-*V-L��������1� ��3�������)��;�|�C*oe[޺���^�5Uc�\��+��J���b���R��r\�� TG�g@#Xe����E[�����)lr�,����=� K��M�j���_W�������b ��(�v|&3���&�,�-����_2�{�v��6�g�b��!��J������^���w�G��*<�Ϥ;�~)�!zd+��HD��^X����t+���v��߫i����@�	E9��������^CoO��p/�g1u�������z���{{XM���c��6
����72�(�Z�k7�S��?#�k��^��\n�3�f��Q^ߩ�b��P�2u�������[x{%��Y֮����d-�4��%(��6ǣ�y�Y⎨F��\�ź���v�#�	z���%�IdF!��P6�m
b=R�޵��t�!fᐘ�b$�&�E��a�\����rAA�	��1;6��}U='�yBӪ���e�͙ǳ��ݒ�?�7�ͮ(S
"���V.q6w���gð�i#������ $�[5Jgv��O��@˃�J����5�k��P��������[I�?m��>����5��Sv�,Z��D�:������i^���r��R�)��_�8n6A�ٜ���&fg��
k�9y>�>�.�c��[�8�q6�!/:�Bܢ�J�˲��:v{�s}$x���$���q$��0�%����cT%!F��PujJKH*O�q��k�2��T���^4'-Җ ��wI)�>|���?��@�v��h�҆�N����8�m�n$u��C^VNY����a��?�zA�_ҳ(�	�C5���ޣ�O\�CZl1n��Q��x͗̂ﴯE��6i�\��3?��E�R ��EQ�>i]��*�RA�ݭ�aO�Y��/��Si2�2L�D��|w����PS�P97Z-����4�;&�c����������X[M�ⷦi(	�f��$�$���'��RG��A4��#�/R�y��_��J�4��0��d�M �''��#Vqi�Q7ї}�A�XlǾ+~�4VEwl)�`v�k�����(��F�[P�c韣qq��Z$��te������loӫԪ �wx0�	H\#}�֎,R���Cs�%Ͳ�*,�Nl�3-�$�0�&��;��n2��rJ���}�@�a<i�r�eu M7�2��X��?t���}DӒ�g5t�
�^�_��x