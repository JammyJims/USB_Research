XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������o��X(G��������P��tx�E��|?f_�6��")����
 �^=)H�4�>� {p��#�2���ʝ�~��k��؋���bn7\Ak'`5�e`�|9�h��Фvv-q���L�&���SBU�I�h�-y�"�v��!y���X��g:P�cڄ�&����LG:w#�>g� }�`c{��0O��D�me�R墫ZS���ǋhu_$���h�̴��q�v�
�� ��̕�x�c����"�<c�X$�a�hkO-�&���������U��{�{p<Cp�g�[0e�<�~��94x���6	9��l��,,��T璦���N6�WJXX~��Nk�{����$���Vo�v�B���S�̟�- ",E%�!6��dD�U�蟀n�����c1�5�4��J!�r;IR��.�����Ƥ+c77I���~}���.�Z�u��T*oB`�o<R�Y@b�@����x(sAS�c�y{�}���mz����0��d�`:���	bB���u�8��hS�^�S�@�_��Fdv��������3_޿��?�Ö��8 �J������D�m��ҽ��0B,��r�f>�q��9�#�L'�����f�,%j`�i����2�qB nyl��l�A]V�HH����Q�c��f3�2PO�����ܷ{�|�*��h���5�����ߴ��g�x�����y�33�x)���Zk����h��F�X��X�s{8�8)���x�sCs4<�D���ۂgc<��Y5ﮈ��$�XlxVHYEB    5339    1450�d"��6��n莈�4d�s��	��s"L,E��e�[PG�=�Bp�E.ީ�(Ő�kY8
h�ͽ�s���ɤ&�3z
�Y*.I�]P>F8#~erE��i�Jbi6����]6��}�B"�2j������C��e.��V�Ҏ���L��rG�$r��q�\9E��A@e�_�����`�C�v���ş��EC �Z���s��"����k��~�̉���7�����h�.皁=�d�Ӵ�i��J$�� *��Ƶ.-|���#�z&�\�����a�PGJ��{B��u��ܛ�+���nE֫�``h��	Nz�9y ��à$E$Fy����w�KBKf�*��h��lȂFtU��(<�!`��oK�h[��~"��C��<H"*,�.���0������o�h=�����.����~�;��U���{ X*�N����$}(Js�5�����[��NA����[�G�uw�u�=XG.�U����%h�@�����0�yq���n5���;����:�[Y}�e��{��׭���7[PevF��f&~i��H-�]�gڢ~�)9�?.���z5�K��)��vqW<�w~.p5Y8;��vޑ�6�q�!��x@���������?��y�*V��r�u�/�r�pX�qG�WY��m�'��5�^i��<��7{��˼���)�Z>F���e˃I�s��'$ʗ���F����J:x,^e���O微\�!ُ��t�}��@������"��P������7��j��ۉ���I:���J#�V�~-���8�{(�G���i&���@��C����(�&�����n�~(�r,��Z�S�~�Bx*�Ȼ���Wԕ�ϝ�0y!g�l��Т�T��p�^�E��?��9)G�^@fk2��>�����-3�[�ko�?��:�С�w�܊V����雯ʗXG�?K��@��9W��h�����u=6��@{x	�˻�t8y9Ξ#�c��m���N�,]NJ�
��!�g2�� y�IA`Ө������Ejzj��9��Y�^�$��XeAP����t�ƪPS����O�D����=�f�Ա���T�s4_���4�DM�n-����C���J(!� J�T��?�0�u.@���k�hb�
xM|��[~�UEuſv�z����i3|AR�+�:�!˺S�efY���"pX�H���69[�-��C$���1�%b*v�`�����,���_B��%iSQ҂ń�mc2�SC���m����ښ���0NQ�>�6�Mn,�2ф����?$Ʉ�_�ͼ��SPj�0S�⍔��cG��k �A.�to0@�v�PD몷�.kt��,F�k��4Z��w#�H0���0s/ml�sTo�	"�+-͚�� C��L��>�(��"J"'i�ic^:E�͚4�N֊�HT�Ij7� �
?w�39�+2a��D^�C�o��`���-t�9��C����6��K��e�������``�KY���d��B������c�'�G�Y�����q��JDL��TN�)t����Œ�Z�yӟ�_���Q���OR�O��I�ˎ��CWW��TdG*�<�b�LP@5��WA����U+*�A�2 F_���9�Bm��Ŗ� Ry�Zn�Ŷ���[O�^�Z�o��O>H��i�D�V�q;|d��i�ї9���݊]9��粍b�\eX�9��v��Y�p�.5y]%�w���Z:7kl�hġ�o�I��G\w�5XF�k�.��p��H'5vN=�T~��8Pk��qKHF8�/�F�\n$�ljv���j�4�����d_�����.7�H�F����2#{��裁4 VoF���Y�˻t�j��f�����{��ay��O�j�F�Ή�sxD����R_�����D���;Ԝ�������Qį�l~�;�L��)j\�^��h��#��5YRN�6�m6I��x{
<�_G6R�Hc�g�*j������X6)^�
]��ѝ�<ɸ�1wa,W9\\J�:�R�����:fU�ٽ��(����c�!Ȳeյa�#?f�ov&����q����
}�B��2���"4�W���I��1"O�wD Q�P�|��Bk�8�Y�GX���x{j6;���&X0b.&�ӱU
�]����i/ ��g�^��Հ�/*��$l��H	�]�O~�Bw��5��a��iҊL���&�3�4����/�CJ�$SʤR��IG>
�\z�?5nU8E�R�B�9�T�]6$��ҽ&x�Gup�:3����:R$T�Զ��)�h"��Q��/o����0<��U_5����J�[5L^��x��6/̜=ma���>a�h�(6�hn��JC^��ڶ#tw����:�~�)B��>Y�����p}�#�U�D*�E*ʰ�ٚά\������0'�a�"~8$)=k+T3|9�k��zOq8ie�*�K=|z��g{�R��k�a������v���+X��8S�k�#B���
y_��8�=�m��܇��=<*��K�T)H� "q�~�Y{k�@Y��N�h������K��ǯH���X�nbI���\�6�����p�ӝZ1']#c�4�&3��`cC���_o��m
�˪Φ�Q36��ܘ��	~�P�i��
l����I[w�;eCv�\pUhU��dveFi���",o?:�/��U�4�1إ·=Vl�Yx�֜![�	^����$�Z��im��ߔ�Cg_������$�@�����Ɩ�n�y}i�y�p�_�$B
����@!��O�����#RX�6� �B��9�吠n��Цmt3����l,���^����?��Ntues��i�����=U��:Fص"��F��R� �t����][4���,Tӎ�g�|x���p�2�αiE�����6W�	��.F�Q$q����W�<���ȏ��Dz��ϙl�xR��,
+���6l>K+0'?�|�<~N^*N' ��&��_� >��(��p�|��My#�kH��i�|W�_#C��*1� =?���B<�+�jLl�.B�q$�~Iuk�3��� �¿[�������c4�ꃟ�]dy'9�̯WFG���N�s�����݉,��^b���Jm9�~8=1����mW���5���^}�o�˧�M����p�(>��$בW����R-:mO�9�-�9�R�H��X�̊4l'�)�j�"��B�}QJ����a��}�ÞE>s���t��9��Cӏٙ��y����E	23�c��.�'�����̘ J�.A(?%{v�0ӵ�Z��]����Ìz�kq͹^���Y5V�+Pô�oo��ʹ���� g�Q/⃿%o�㨋<��Q���;H�������.T���lk�y+Y�&��-�ԥ��2[QîcA+�2�Tէ�#^)])�0'�����Y�c�	4<�Y�O|�GEP�+չ�PD�vM/�mГ�?(��U$++���@S�3����,���|e�� 8x�dw��;ω���y���4_�h� ��
J�*X[D�%�{��Y"�{f_M$:A>i�?���i����I \����L�6�0���Y]�ϧ��2��^H(T�E�2���5FF�F����H[��F�<��bɈ��9(����Ѿ�v���R������������Ղq��Gȃ*A,���BTE�I�Ū+h��a0)r:)�ҝy�W|�
�KQ���2��e���\@d˫���--�k��#�LtG{��N
��E��_h�բK�Ҿ!�V<,d ^�
C�""�\{UA��
b<W��8�jU�~�q��
(M���@�e"�ޚ^[eltF� [ �o��>!���Y����cX%�J@$�n�ʰͧ^��6�֗�\+�M��ꉅ����|{���\E�L��<���'4>�%K,�RC�-����cH�lHԵ0�)���5� � �P�▎�rǬ�+�zQH5��jѻ��Ĝ�{<|>$k��>e��$����?����)�|&#���z/d����f��j�4J �g�v=���C	4\�*�,�S�@�K
�^x\�����k A�K�H#�d����Ȃ5z�B�[`�/�C��92u�9�/'���Ȇ"~���W�˅j��F@� _'^_�B!�r��=ht�ƃ0�yA�X+iv~�A.�N�v�<s=���8�����Q��4b�L'k���G�QY�C��2�V۠�9���6�N��Y���5�<���v���`}-��yGm�^S~��l�CO�C2������U�J-��t�C�^�"˦g�L��v.�W�;1D��͹�U;ĈEc���$J��#P��ة	XNVQ�mV�ˀ�:�Z->DN���0��lu����\h7}�x���u�9��nHu�w���~��X5x����8��|m ��������Z�<��{x����O��ȳ�q�a��̈�tѽ	I�qh?�	��"�i�l��g�6�PI���/����N;���a�}����Vj�&�psԚW]f鳾�R*YC�&T�
%�	�̙ҟ5�;V.k�ɺdV� h��/>�yl��yD�4�@҄��|z?Xz,���o.��"��@�e�Q�aE�3�J�S��CQ t�/�|9ȡ�\h��BMC���D��1�YH�T�t���ᶷ�'gFХ���>�j$���4�� *|��$� ���������ߡ����V,�~�Y�eI���|���i&���&s��1W�G��{�
�Y]P�(���:g�T����`��W��I�d��h����i�өF?s��(ۜ�t�kw:(c�n(�#������R� kì@� ��&bW�	 ʏ�*���) �a�	{JjD����-�8H+��̪\���ٰ����):Q�g&�;�IXj��=�]�i���:Ɠx���Ns��M5:�;�N��#q �נ^���8ؽc/�:�?Fʜ+��ttH��'��A���L�D��,z^�M�Z�� t�P^x�u�5���T&+ ���Q��+8b,���~~T:�V�i	8�7�^+'~���^q�I'��x=���L��ٝ�V/�hA�N:� ���xI����U������oև���&�Z)���sN�d@�7ѢQ�Pm_Q��r$sȧJ�