XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J�-�d��zO��&@�Nǥ�ꏅ8�z�u�vy��r#��굮׎�B5�z[&u������1	�v���V�#{Ź�}�s�!]�'��0�]�ߎtW������-&�~\g �hP��і�K�!����MD�j��[�pb�a�����k�ɊA�~�ܡ�%1\_\��M�f��y��ฆ#���W7JÒ:5��%0
�i!���#*ĪÍ��[�`q&��J�D���\�v;D�Oh�&X���T��/�`�L�ޱ͗�����eQ���_ʃ%�q�������~�������r�d?�(�����5�~���Yһ77��H�z���1H�pk q.��E*	�,+�,���MP(~K��ljp���Éq�h88I��\��:�+�$��@Evo��s����
���m7���Z)����aZ:<���1u�w�Q<e�M�ssQS��4ѝ<ݑ-�5��挱���.��V�`皦�ی,�q����:0P<��-EO�r:4�����׈�s���������"T��JcB�|n��©w1��u�����Tc��#�;&�p�x!����/�Z���!�]Լ�9���pt!�_Z���qQf�ҫ�譃���,�$u�1R�a��O���?`���9<b)c�3�Y�q}�p�R��zvy��:
���e�V��X�k���Qk�a+�4�S�%c��mZ59C�T�i$�$�ǟv��,OK$.P�����?|(T�E֭+�}7�\�l��>9BN��bXlxVHYEB    7310    16a0�C����ҫ/������a�
�ƒb��p�]VrRl��l�4v�'.kF^ ։�u�]F�OT5�q!ݳC��
t-rU�'�.���prNݼ�eW	���Oq���'4�}M�lav����9�u����U�:Z�vY��H�O�e�QX[N�x4N��\�ó�YFN�x:ʲ�V�{��vm�1�j��n^/�u�YFO*�m�_9u���7�}r�G��k�l���7�d�{݆J&�uo$��F�V���
sb�ۣL<Cn�.&�=��eTI2i~q�"h�B��������/���&��w]mGT1��B���3�Z}y���x�^����-H�s�nR�/ͬñպ�K�/�<ȯ�q$f�����qZg�;f�F�~_B�3>��v�R�[��T}ue�|n}�7f�w/:�����j���g{�Ykd_B��}y����z�p�1�M����i;�lJ��a�r��1U�鱮gw�P8���oQ�
����~� �Z� 3��e&LҾ�\����N)��fOc-�õ��qA�-�*��&�!� 8n���:O].m��I�!�����(��� ��!�*�q۝r;9^���K( >��u��,��)�P���O�{Ѱ���u��Qw2�`�9X�t���� +i�����48�_�{k۫i>��\�/�(��#�\�$`���eR<[�}���63qal�����t��8?��,����v��S�h���2m,�����*ʟ< �d:�����<}�*�-����pV���ɦ^vT6▿�{����?M@��GNÞ�>J8��2������:���A���|TV�����
�]'V����q����W���!�"�	��V���!��tΨ���L��(073�;g���yw e�ک���~��1�ϟ)�KS
M�e�Ip@��iɐ��VI�''�����aHƽ���zW��,��Xh�Qo#��ծ��7ԣ�}d���e���8^�ªHj�`eH�����UƤ�hb��I2*^�Y0HX%�� ʬS��*�!�����
�j�� A���#��v�\܍Åz�HZ��d�*hRu.���g1����r�\y\a��J&m�
��գ�_������.�b��^1�egu�1�V��u�}�߈�����\�y@��D�������9���fP�Ar�	o5Hu�o��/~v�Z^ü�?F���Q� �]j�l�C"8�/�{��})R��~�;U:���`Z%R�����l�C�;G��{�k��Kx� u��=�g���j�*�2ڷt}V���>�y,mk�7�X�6�����X�7к$����dÀ�� ~E;�Y�9|-����%��6\�q��"���?����J�nւ��E�y������(��4l�`�'���|���_�1;�5��;3���:�#��^fAtq�� 4�Ǧ�%?܋A��ȵ��)����1G9���ҹ��e^�?��n��-'T�Ay�ԇ\��ǌ��UZ����h�y���F��
���-sL9�c�D̗�س�0�{o�и�Db���p8�Ӄ�U�'��4�:g�ř���f.�4c�$"rᠣu��U?a�Xvy-~L�-��.`uፉU.�,��B�1;���x�N�Ԓ%4f"��u��7D�Y@:!N�<����f+�?8"���z^�U̪܇	�` _���_k�H-�b柔��������sMdh������OK<`��ff�DH�p1o|�������6`D��Cq�B�>Ъ���%o$=����*�z��E�NK;K^eQVʛB禰�7<q�g��.~e�42N4���S]{n�� �X�y���3\��Sf����*S��T���(s�\i'�FU�����Ǜ��b
�{���A�*�cMd x��A1Sfa��כo��`E~j��ЁR=�}��uP��bS��j��p�vY�x-� ���2���B����ڃ��\��Q������RRu>2�!�1\�>3�K��5蓖��Śc��!޷���6oO��!��g�=>�BW��Ӿ����bV������TX��a���I�1��q`ICHGD������,�n��|�޳���b!R"�O8�؁\�#H����*,��{fNE
d�b��"3k��k�_:�'���~�Ch���"�X�yAП�̨��{)�b�Y�i��X��� ��B,5���q�0��H�ʪl(Ʋt�Q�a 6g8anK�����k1���d�Ӈ�i a;AjyL��e�@{���ZH�}QZ�ΐ����_綰1�_	a��Fc{ /�=����YtV �Q������ ��Q&�7�t�+�{�g��G���s�0��|�y�.`�Nq� E-��ff�ݜ>]���rD��1t�k2������?Ҍ|�$#��4��ȓ���y�+,b;�1Jt��eq�6M?�vU	Ɣ7|P%�*GA��%�Jx�ҳ�IMi�mS�~�2��TP�e%�#�!��v8��o����LǸą��P�0�Cz��Q
{_c��$�L)<"ɞ�~����麷�ya��(���ʽ���7�ʍ@,�E�8�B}<o���/���;_殞1�GF���$�BU*��M<�T����xH��xPi�)V���i�����	v� ){�H���3Q�Q���N��'5G|��[n9��ϝ`B�F�����c(��j��i�v��t�e���!GRF�ExKt�Ups�@��Y�d�]���� ��I��^� �Y�D��D:h5�n�yT7��R�C��r�R�Y�![b��/�NK"��p���o'?��W`�z�X�l�hr���$:?��2�	uNw:�n+sJ�7���n�k�i���Hض�	�駀f$�.j��.0�sJP��xǳ1������k�sC� �7�&��{&�`���p��8'�~S�����eq>�ￊ/^2���̠��<�۩�8�em�0���޲�.y��X8t���,R��%�c��	L�-�Q�n�5y��A��Lt1|uCHc��ӷ ?#$���p��2?������������)��o�T_L\� "�����[O�K{^٥ݟ��_	�Μ�bo���e���M�?���oY�"4�"e�����`��ݧ�Q�}��ڙ "��9N�Vb��A%����C�g��ￅ���j�
咨pݲ�)�+{�P\h�s��Az�ǖ@ܚ�HHO���ew��N+Pا����˹��w/�������� �| ��^3Kd��Pr����b�	��\�z �	���؂��I��{x�����5��Qӡ���A4�
�NS'i7��vF8yO�I\[�;�3�N�Ĥ��m��񛽄RrJPR��ɾm=��XIO�U���	`5���7f�5<k����@��)>fȮյ.�?|P�(V�.��5�9Ӱ��u	����J��%�&�U șl68��l,O���<gĲ+��l�+�]�����PŇ��h)7��Kp��v\�Ld�:�&[��!ROXUQT|�h�[�W��4�⯙k�|J,V帎�FY�����>u�[���r����,J���m�Xpw;8:6�M`Tm�C�|B��?���׸1�$�K�<��0+eN�~O����_�v�f��::|�Ux?pIR�X��:7z���5Q(�k�����vC���M"~�X���N��K�/��I��?��e��o׋����܇,����)k��~�~cm(�X��"`<E�'\��cass�F-��S����a1Ï�q[�=�14���s��I�Ƚb5��G�^n# Y�}X��b�������6.3Z�@���j@��8G�u��!_%`Y�a=�8Q��qC��:���c�'T����K�������~�ٞc�1^�
ECMt��8}ʺC��N	B#J>����gZ���5oA�%c.0@�MN�xW���v������G�N�j�>~Fl����i��v A+g{�X��$��&�[<�g��S�%UO�v�z���	���ZY3�>��z �ѫ��#�/����A��1X�~+�3Qa���'Ha�4c�őp	��ԯ����r#6^�e�}�T��&�D���^�㡫_�/����Ik��H=tW�og_(���j�_�G�W�!�l����#��t(o���Z�*��G9��W���Q��f�T�2?�+�,ǆ��Mڬ��,�%swB��ǣ�d����Vc�j<�7���Z�i�;��M7F��9P+5���D5��]a9�j�.a��?�t���@k�]�}`��}jw椱�	�����\���_���3�FKF^���!۾��Կcoec:a���2
��i��&�>Yab��9��x��������_+�D50�`���3_����1>�A&�%@5mB����G;={~d�3#'�WHF�]���XA�-��צ�� ���hXNz�A7{�TOH�p6M.�M��P�U��q5#�>l�Au5R��Ňܽ�{��>Q�ZHw{4�.`��l�h����e�|��+�˘�}�|Tڕ�\�IŌ�)�B%�[�f��ߖ@Sju����\ٺ4��^��4"6�ۙU�t�6�N��c��B�x�+@:����*X�p��rYxA��v�t�|�2���3���{.�~������]Mp��ī�{����W�����Cۄ�˯/���8	OW(�Hm��Edq���;�bm����W�-~���n;5��\���4F$^����r���4!8�.�t�O�u�����s�߫ne�t��	ޑfꗓcBN�9t+x~X_��\ѓm/m∘^���v���O�(�:��B�K�q����E�ы����x����8B҂hܷ�o���ű�G$�����˦Q͢��6�K�S����'e�:��3΀�id�Ђ�4�+h��$������2� �z9�����5���.[Dc�ΖHJ7�b�������=�.b�W2�
y�t�Q[(�r�:�;�5F"{>�@A�x&�#���sM���Ԛ�ƶ=�U�%�S���p<K̢������I�ƶ|w�:��y
����{|2M ن:�tx�� ��s7�{Ii:��[p7~כ���w %;�� :�|�N3Jd����5�����Ѵ�"�㬶����`0���
��A�]n	9�t������C��+�u����г��*32?�����.�"��s�2���p���X<Z4s�NS�'���a�]��Y�	�<0� ��T�i�_YY�Ĥ37�.�*��G�Va��2��=[�G��� ���?�D>l�u{z�l�DM51�X�C�Y7ڱ�~����U�诟R�I��� s*,>�EL��H��s�o�S<�e�?�}6�e�sݦ���~�ҩu��t@L���h�r۟H|�P���Ic l�kl��rL�m�hn߃��B�V �zq�Ī{�Y�D�&)hL@���S0|�7I��oC�Xj��Qn�V��_H�m�O@p��vJ���3��Yyd��_ꀜP^5��*u�y��:P���Q\���<\��Ιc�+v�߻0cK������"�$;va�Pդ���n[�� ��τ7�_*xj�s�j�a�c���w���{�������Α����{��/��|D��˂�PZ �k�tO�-�yxʾ"b�G9��	^O�ݗ������v��v��ZWL�f��ǰ��!ܮ-ڢ�[�x��e��	� `��m��,Ć�����Q41�-���