XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~�CUT�q=�Qֿ~\��i�lY�P웜��ʺ�S�������G>x���i��?ջɝ�3Zx0�;��Tp�/`B{"�쩾�TK��;��8_=U�i-���!�߼&I0����e�u�nGn���&˛l
'C��t�`���`V��Ɲ���6�q�	+�m��*iPa�Ǎ���v7EM�B;�$}m�4��~^��B�"�C𮿹kk\��Qᳫ*@yע�ZCz:DKȨ�ցb{/q||=��^���E*D�O��+�(�N>�q���"��{�ѻ�%5�%�>�+�D�:��0�7�"{
�3k�(�˭=��W$�	��_�V|�
��i�N�ݬ���'W��J�b��?�`
�� A�^�@�������V4!�k�D��Lg+)���˕��X� |R	4�a��`���C�4;�*�qx<l��T��|��עh�Z��~(���C���MȢ*:�ѵ�D����?
�,��.z�7�&����7!I�§��(���n� �g��^>RMRc�3!�W�wP!��TORB(�<�W�\u��-Y^v|}��{B�/��?�؟^��c���
���e4���P�0ѪP�)s�W�(�4�YF�\1�}rK����L@��x��06���$0�A�W��; ��Ӛlدd���Wp���g��C�t�>dz.�<�B>bj����яM.��^��3�����g�Έܱ������� Hg�L��mڈ}iFH�Uy�A����*^y*<�XlxVHYEB    2230     9f0�\���%]�Jŉ�!��Z<��vO7c����C�5�D�7�Xh�u�:��8]�T|B�e����]�TC�Qt�3q�(�+%<�R��J		�=xIĸ���L���mF�ck0J�'�7�ogW�R�߆Lg^��m[J�$�W��yDi���7kJ�!;�B��[�O��z���o]'{�[�ٖ%hU0*��>Ja�����j{. &��L�������ߛ�U���X�wN����b&�*���Vt$�$Ϛ��������f�P�dZ��aJ�)�tZ�/ �����n�O(Rs�O��S�����[c+C�FnR9����Fik�jiE���5rD���k����Y��_f�,�q�f��1^i;�͏�D��v�pS�u}���{v�3T<�A�wƚKx���e���=8�]˝}�+M���6gO�H�t�����Z0�-6�WOg*���i��
G�O�m[�h����� �ܷ-�
������D��A�]�����.��\MG���ԋ�ҡ�KR��D��lKm|��$���|��ӡ!�^Ts}�'�MQ�S���8n�'+B�NO=3�_˾!���'� Pr�3ە�9C�����*�G��^�e����鲞��Z�J���7C�54*k!��n���:��a��ZT]^���_��� �9����]g�s�A�nqy*���$�K�d�3z����4$�J�*W�+����q~6���Sz=~h���P�:Hߋ 99�&"�������5�7�ʹ�Jo�����Wy�ǒ|7k�f"��:���6y�,��WE{7v��h�MRݺ;v���9á@9c��r�U�����z�n+k
������˟m��,������$p��d�H�E�"�ɇ%i6�,���R-�S~ۉ����'�}��_�έܒ�%'6���j$���4yxO�g��r�n\��xֺ MЕ��]ī��"h9�'�����LC�0�j�x�4K��%g,�+Dȩ�<�M=�$�x��Fd��]])�ǣ��"5k̘)�Pl�`:m�P�%�VlFna���t鎈��)|��@y���q�V&g?�IZ|���6�N8	�s���:�1=%嚚+fe���St��y��eͽ*-�����g��6��d�eA�W�gV'J["����A��LF�l
ƻ������"�����,�U��nɉ+�ݷ<l��P���9FoP�z%�޻��j��QC�:�WZ
8@������:OQ�Mկ(�#�x�bCH�s�D��ݡ�綐	 g�<,������[�?:�;P��Ǝ9N�:�K��+ܔG�M���,�TÂCO+x5PB.{Ў�Ufx�>刃j'�`$��V��흠kM�IINqYI�w�1]��Z�EC��{�^���.zeU���#���M$6��~�X�j�3.�f�p��ϩ�'^�X�(�8P���~._`w�lM��~��3P�aٱi L@����Ւ7����J���b����������ݎ��b��E������G��
9p�i
{��=>�H������������3�$��ܫV8��$����ё.��:�[<���>Y��@��Í�"�K��fw
1覝�����h_VU䧯|\�0P�{�畮$���Ȃ\��w)������lvt1�P���<6�V����0̕@������$���J*���/�����_)֫[� u���c���C�:�F`�ҶatW)I�H䀫��7���MF�����b+E@��~���}*��Kڡf��\��b9�"�ͯ©-x���rڑ;X�I��N���}'
�z��\�E�[+��G��_"�丼�����nB���J\���)Xh�=��AE�!1�!c��G|��v��:$�L��ȩm�����}i���	qe�|���.�|s�w'���o?�*T�>���'���	�U4P��ȂN���a}�B2�y+ ��G_�Jlx���X��z ?����J� NE*
�_x���mANM!�a����!@�U� ���n
��[�Tdr�+_�׍MP)������kd���a�T�����	�up+4W���7�ݖ}M�U��gZ��垇�~��#'�����6B�E9�A���'G�z�X��w�kA�s=����	H,Ӕ���s��:�<g�l��>��0/M���_��x�t>)��U�����0HZ�X( � ��*{�_���g��	jї�O����j�Q5s������W��%T�82�ס��]��q�$� �q��[�z/���{�'�AЮ׳���Ci����M�Ҫ���6/��r�Q+M�,�O���
H�U(8[���J�=_��_zQc!�݆H�G0��d>X���Y2�}�]��}���ֹj�f���per�,�I�
T�PXV�]�w�D2���R�#��	L����x�K&<��U=R��G�M�pF;�i���7���T>p��u�JO�j�;�{Jv��t]V�C�-h�QN~�G,�
9�