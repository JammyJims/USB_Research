XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�������r~Y�(Hy	���K=�ϧ��D��H�ñ����|��=�1͈H��!�@З�k�:��I�c��F���R���47Y=�&J��%��a�R6�啲�����#;����I��Ͻ+̩ň?�c�9� �n��ܠ�p�)	Ȗ��vi��o���JO4�һZ�+~s�&��`���w�Ҹ�zqH�"|��k�}���j��� Nz+��*�"��,+Y�e4ETU6��@z�p�'���s�UVjk0d��}	�T)⥃��ݤ	?.RkT	���t� �Ͽ�3�E�O��)B�;����L��,z�
��|�Y	n�c�DhL�8\���k_coc�v��C@H*�\�M7U�)K�,Bp��#��A���H��g�g��=d���a�n�ʝ \�uB8j2�'�N��:s��|����l��3�P�C��=�'s `���{��-I7
��� E��#�>F��os�}�#@��$�5L=�n4����������O0�s�� �]��K��p���#��0A!���F�AV#|�F�&�6��ѵ��Y�%���K}�
�hg�x�5f��ϖ��OV�e8��u���ڤ�jcp����@}/�(��x q�����4�c'왋������DH��
1v� ��Ț�e�:ͽ��G�@#s4����D�=$=� n+���Kw�H�e����	��vh����W�/��;n!j��7Q�8�;Г��~�u7$.����hqy�Կ��-Py�E_�Uݴ�A�Z'��XXlxVHYEB    43ff     d80y�������c"�o�6�x��z�E�\�r�-�m���)�\������h����^3dfT�Pm���_�U
�>v���S��rhI�l���8Z;�&�{��~j��J/���ѓV܇�����}]��ST���j>w�^�r v|���<[����E�lٕ�r$��l	�s�S>V�cUF�4�C�6�e��G�P�-�#�FO�����#x�|%{�޾�>��( �,�:�8ˆ���S{��h���~nL;�s�	u���?d� <i��P�B�]��	�W��oJ�x�M��lB��Cp'�։w�9�HΝk�L*�Ր�����h��gk$������p�*tyu�޴�}� �~��.����# J�e<����lׄm��){p�+۬�μ�entI���	��]���{Ȓ�mA���Jq�,6��|s������o�-��D�gJT�W
x��C�s�ʝ@�D�a,��jʎ=qk�ǻQqYJ]Vj0\_=:a-�&�<�&8���"���2c�Sy�����\֭��9�c��ow��)�3��t��$I���j �9 I��e�ýU���!�i6N5iPd|�W&�!4���+
�kα��7��N��������>h��dk����������W�` �݂�X��+|�����N\ŠW�_�O��!-]_�����Q̙�D�W���w����7Կ@%2�A�	����L�J��i�J,�.���y-�vM
1"�}�d���oĦ�������������sy����۩	sU	�#�.3& ^	��9\%гkw��I����a�\��Zx��Tkj��V.���ol�Y��^ �&f6�P��|���:�y2R\x. ^�pcd����%F�;�99��'��|C!();tP5&��b�������
��j��G�'�+Yaޫ�:�]�� �3��" 0��b��<���"z�(þ���~N�Sc�FZQY" G� +ʵ��!�=����Z��O+��d�/V&�bL�S��4N�(��3��B]>��7I.�����	��ݤ-I��R%��tՈ)x3n��-�.*r��I��+Ke�y�65@��8�M�ڷ�u�`v�\/��KSW0��*�U�
иb7���+��w��Րd}���O�^�D&e�2��Ѓ�ؽqH��*�c\���wG� �.��v�`O�6��w��9#�@�nl0��85;��"<"�7��{��%�T�Z��><!� JHd�3�xk�G��V�V(����i��w4_1�,r�LS�!z���-KX ]�����K����T#!<m��j�{E���"�� }��! ��V̓d�[��x�{�8�����e�=���T���|d;e�D�t�2�[g����C�Y3w�O> �e)���U|�o���'{��O�Z���ʃ�*A�GH[�s�3��E�����֟��Dp�Oy��h�7�O9e$�m ����2O�7��P�G�X+;�LYW-���qqՉ�c�錿6���P��J<&�8߂��W�5E�z�\��vM>�wy�qN�Lw"+����r4�����M�t� [6	H1y��'c���;j�T�K�z̑w�6�a�&t�Z�X�G�4�ηwƅ)H>��O27ULf�+1f���R�髏篦+�{��5���U4�J���U֋P�9i���7��C��ถS�ڨbw�c#[����<Ń��Θ�Wz�.��o��v�IL��"kn��Ӯ�i����8�F�`����z���|�Ԝ���f��2��O,� 7mFgYl-��8@"�kH�7�.='����xY��o�`,�u�P<ƈ��M������4\Lϼ��ي�
0[��Tn�޼cW�PkC`H��I.!J���y���E���P[��Oh�m˕c+[Ҩ��ا��|/ڤ�q3tU����|��XuA�5�z��6e�Kn✵��n��$N�EG9�[�S���0rh���5�fMđXo18pF$f]��p&���sˎ��Y�ӆꝈ��oἏ��<���.r�(��z>�E��´���O�Vׯy�jX���׽��2��V����?��P���2�;�§�U����k�RW#(�FaX�_�w�~�=��E����?n�����ۀ)��M�T��٭��+�WbJm�P�}ؐ����k�7z���\�][�KiSG�d�{֗�LhL�j(}��H�fO�ևߺ���*�g�8K�#�6���Z+���r܎���c��n��P>J��z,|�I@r`#Q������KTD�[63d���"1�F;9�����R�N�^����A��P#t�FS�u�����UT"�y��������k4��.�+���+��Ot"��ʎ�Ql��i�B�&E~�i
q��M��=��
]S��y�Z��CR��b�.�c"ۄ���t�x���\\4TsfGC!3m㈜�w����>�8��_�[(�������-��(�/4ά̆]���ǔG�P����1��Ϛl�h��V&�d��|�l��rJ��4��E����
WoH����ޟ1��SAGňʉ����c,��_ܪ]�me��PX%�5B�!	H���S0^��fw@mH�J��:����*���"1��TG�m�VEYr�+/�̒\PI���
��զGs�S���[t6dȿۿ�D�؈^�4����|��âS�y�ژ���K���0��6"��-
��9��i�OO��@r%mHNm����h�8R9�-�����#7���n���Ooe�Ψu�X��H�_��Qo_���s�J� �|�YrGՍK��=9�p��Оb��׉��^��'"�[�5���ݕ\-��M��cpLM��f�k��u��e�nU'_�O�WX��Az��8}#=���D"�͊��ے�/Ǳ>$���XO��B�-��q� q����R���_ptG#^2Cy���/�r�5��F�,���k���%�ɪ}��9�xx^q��<Ǝt���{�hI8T#� c˻/�=� �2����!٩�"�*_6k�uۺ��'�� R�Z�����p��nH٦��oYD�:����n�.+%x�����ɷ�P����+��O$��O8]IG�����tib! �gӽG���U	ʯݦ�Zw���`�6 �ʋCX`:��'w��4�H(�V���,�ESjO�%�|+t��V���V#\��'V�u�*j��Cx�o"6*0�Q�3����;P?EKZv���ۭ[/�Ul���ߥQइ�o$���V��W:���0J�+����|~Z�0��.�p��<��\Ig-��F֩%c�;�+�v(���m�H���z)�o�y�QŊ,��M6F�83����,[�L�B�b�����A0|��E�������8�������6�#ɺ�