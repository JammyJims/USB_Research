XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���l����-ju��h���	J&B��=�ZEO�*w�����;cS�D�C�zWm���$4ٕf��I˶����h�,�9��\��E���حBX��-;�	�N6�'I���_)��q�V�{{	�N)w�1>V&i#���#�hd��"5����#������!k���h�V�����JN_<aN����Э��Қo��oP䳚p�15ҁf�h���[�4ш�J��~^�̤���9f�Pp��BДU�V������JF�����)�m��4!b�����~��w�^L�׳�V�"N��a{Y��h���'��is6�158=<����C�}�׹i:� �Ox�n놶V�����-��`s�'�e�$�2�@8)M.���u�Lc��TnA	�ZP�����J�vM� �`b�2���X֖��B��@aD���O��-?���傗�7
s������É�A���wb�{R����S dvf�V?�Q�g-矡,g��W���d��6�a
W�bETz�e,D虎%9z�VJH��t�5���9еQ����2 �1�uVr�H�D��p������=tEyu\��d���2���x�S�Ä��_+�L(�`	DYN��9�ع�gZ�v�+���"C�<��E�=F�^�5�2�;bz<W��f:��xS):ʉ7�G ��ˉ��G)�=�[��?�1�$Oj�׫���/��\�O� w�avv�y�W��֐Å����N�b�)N��A����+��54�H��#LE�!&��TUXlxVHYEB    fa00    1a0061b�:YF����k*�u���LK���S;d��apБ{����eAf�S����_����bnl#��*����'���-T
�]����zŧpX��R�����`K���*��n$B�&::�	=�/�P�ߙ�8��:����G9�����|��ũO\i�0�y.��gn�d[0Iz�@{��Ϥ+G�좵��l���p��~���p'K�M�o��euv�O3�A���P$���+i\ʡ�A�$���;���o��Hib�����Ԣ�sV��;���ֈ}��5�D+��#�#�7�`�d8hE���8o��-i(��ؤ���.{]r���{,2R�;�#��`�{�EL^�)�y�B��� ^�C+���J�����`�\�J��n@b*Ϥ�|�4�M��'����@�r�2�ZI��8Ns�V�՟vz�w�|���p�6O��y����C`l$��:R6E����8�SY��lo\���=��j�Gނ��,�eZAxWoN� $���b�6�?��nq��,SNulv�i� �٦�	�͘��llV$�Iݳ���/~QQ9��@��-�"��4ϙ��Io�Y��w�:D`Ė�`X�qp2/g���q'����;���$�&x�楸]��ƣ�?���a��ax���Sl���C_�)Yw'�U�d��#)���Ӗz����X)h���޹7��r���2�������V3���4�plЛ:A������������Yo<}=��7� �+� qqBu�~���,�������G�f���ِ�� �rq�D]�+q�>Xw��~�ȀKcz�ׂ`#�kEz�K���j�b����/��:��3g,���ej����(r_��(J�I�V�}��Y7J��Z�����0E ^�4į��^���������Ɨ ����'��>�iAz���'h�ߋ�ߦax���#;�ٸ_ZP��H��E�'�b�m�W��� \���t���G%��F��>P�w�=v���C��v���q���C�[�Pp5uC��A`���j�3��U�&Z���l�1 9	�F�?��5�BBR���[�T^�ex6,���"Ҋ5�5-9C7��`����l��]����V*|���H���\��s���	���|�(ٴ�X8{����a;2[���a��_�a!�SvV�8
̑�^���B=�j(�u}�_�n��mn-�ѕ�&��;����*�ku�����w����M�F����0�)��")�!�Hl���l���uU`Pԣ��eq�z'�R^��e����S�F�#��CD�l�H�J���&�n:�;��V[�I���z��xa�P�댫E�|GJ���-��del L�Ҕmp�4�k@�fEGw�h`�b,�!,Dq�����jx���H���_Z�{����u�L�� �ݐ�-`\U�I�]��j}37Ty5�@��"��ǃ�[K�+��Sӧ�ga�������Φ�ZEvзN^�*�M�)K�Q3{�������X�ofL�>�g&țG�n��y+h��V�rl�%�gq'�n� ��t�>�aê�"U-oM�60f�{d'�S�u9�Y l�:�d���K�G`��F@�mΣ�[�0��s8�]���F�k��&4��?��6�,H�
�/58V>l�d_��s?�#�|�9S�6f�B_�ǻ��gi�A�g�XX� <M��S�zs�mL=���<K�H�a��̼h���.J�
% �Ѿją[hAc��@��T��r����@������e�2���T�b ��h6��ѧ'&��g�T�iXr"�I�i��l���N�hx�\ݕ5X̕�����@�zC-G@�:t��_ra��<t!݄�(�������n�b��OE['�ܿq��sf�,��+�'�W�+�gzd?����I�S���"I��s_o��+���?07Mm�Ơܤ.�����cM_����9�}���t	��=��i ZcG��2V�� ���6^A����E��Ro�?�n0�j�~u��{X�����Q�Z&�;�j�q�{R0\��x�
��6�Zf�"Z����bi����;p��#\�'Ɓ��+,υ��.#䣍�$[QK������ܸ���x�@���I����*X�A+b(e���4�g���&��A?�i�;��a���=���.�����1:&��f�����:�ɣ��h�mZ���a�Y$~2V~f��z�cBh{zF���y���q4n9)�%Ҷ������޸d�oC��O����s�ѶN���L"�;ɝ��Y�i�����S�(e*����nl���^��v�+pq��sʶn2�
��k����|6BE�V4�g�:X�0���KeBm�����Orc��Aњ2�Όe4I�0~\bj��R���~�߆��z�G�	�q�+ ��~���pK�̐ыi;2e�
�a�Ǳ�v��z�P1OCT�$0ү�`�i�w��ܽ}��$�bq������.��	�bo�o�pri�t�|��Z�p��=3ˢ
��)����|�|_)��d�s���r3��V���8�z����	7�[�-q ,B�g�]�&�_��\g�Usd�^ͧ�_}F�vj��� ����]��Dk�?��j�}m#-R ���Ѐh?T��ʑRnC�g1���@0k0���_S�sԁ���G=����D�O�'wt�n�,���4��d�`��F�z�.�4=��c� �LeFy��̵��Kj_�����]���A��٘�,vǇ����R�ƌ���h/U�� ҇���^� 2dI�cP��N�i��'|GUÊF��`H^�8�X���mO�-1KJb�p�u2{�l�'�5��㜬k�w� �
�RL��6�iO��+�2KF�)M��@'��O�t,�[҇iF_���=��Rt^��>���FH��vw�sv�ʩ@���.#�h�ֽ�`G��Vݑ.��E�QZ(��d!q�Q��H֯��@��'ri��݆�*B�s!�Mz3`���ۮ��:��ŝ7N������8g�R�
,���g#_���xN˾.N�{� ��T�u���ʋF�HCdöoA<Vh�6"�\�(��}�KG�Q���*U(c�#Ѱ⺝�=e�X����~XG���m��^���cQT�l������5>jk�+3ep�}��!�b9
DWj4�$�/�.�!�]�=k�� ����j���2�"qWA
�ձaϓ�%�j���{WNz�`�&;?'���Ê�vr��Rf=R؝㉰�=��,����+l�ch�Ӏ�I����z�-�)���joX��A85�M^Z�uʢ߄%�Afd��f�|Ȅ~�l^o�_�KF�Tv�L��@��RxmN�'�v;e"�-� k/�|���t��x��G���� ���NuY�]�Ud�ř0M�?�)R���K���&N�����9�X�.U�ыB?%�s���+�-�|IB�G�J��^X(5������B���N�Sn�4+��a��%�=��� Ii��,lo�|%�������)K˺��}�(�q�({��\�Υ�/|o�Wb��m�d�P�ZW�����z�'���Y�ۢ��*���ßFC��LH�9p ���VU�n8��l�.{���-�����K�z��ؾ_#�:��9~6�������+ul�&�
�<�!�|���j��e!*D�*{}���Ӑ��>�A����m��������m���Sv��9�}����wWG���u�G��T��0��ױ�?P���M�0������\��.:�1�0m[,�-�w�j��_.?� ~=��H�c�o�1Z}�KX�1c�t��1׻2\FXRh�ļwG5�3���'�U�D��l�`�J�|&���*j��j5�K0:�R�DĎs��ѝ��0�:{�,�p5_L�K�;�Ƞk��A�t>���V�gb�����)CO���o����y�D�o�Z\��й}�NO��ҵ��F[�ۼ��в���wt �1A�qE����r9������#�-�� �37�,B_��WX����սX���[���[8�\�K�������rX:Be���,��N�P;�b��B�;�*$`f�!���Lt7Sͯ�s
r
'��/~�hu��ɩ�I
�g�}�e��k�����+fB8���~��xAĂ��<xsId���X�����/�#�\�s.����t~� �9�g�k7m\���N����dMn��ܬA�Pe�y]�fA~0�O��1Q>���):S��@Z�h�k=��J �ٲG����#u�	H�?��2�SԀz	�a�����9�>ԜPQ_���7U�/�������,�	��I~#6�]Z�gXA�� �d�tz%1��x���'ׯ�O��*D�޼�IiF4�8�4�MGZ��4Ҝ{�L�h�#So�8��� yH+<�`�g.R�4�_>X���u�(ۘ������1����eA�7벛��Y���N�*��n������lE�s<O�jUo��8�7,̊+����������(�x�Q�2Ⱦ�G��	���ay/�<"����&맜�_������k��=�o�N�HJj�nD�0�4UDrKy̬���1h͗�ƛB�<�ZԼ�A�K��"��RX���e6��\V�B1&7���Ra!8;Y_Z�Rz[-����PE8�E5|���K�3�dH�o�L��bQt�e�{5MHA�3�NX�Bk�h8K��7}Z��M�y�Y��rܖ�'heȳ�∲�����5�xQ���W[�������_� #Qu��.����z����E�ƀuϱI�뽦u��'�ztU����8��e���V�������P\rGSh����ߐ�n��O ��
�~{�$��&�BNi��u�����p�W���.r��	
��+k��S�F�cJ f0���CM�3&�{ڴ��h-�̅�߂�z��n����?��龃�	�2y��ƚ�#>�+Ȃn�Ndf]����zG[�7
��"*_&�C��1�7��ݙ��N@��
n�x���T��ӯSa��'���h;�G�8��\�t,�ăF&���<̆�[ņ��h7�֕��E�G�H��o�)�筋ƨ ��h�H�����럆�9��}��5JV�O��w�G#��SZ*�펻^��`^��u�E�y]ܐ��M����?�8�ߟR�_�-m����KxCh����zh��!5�v��1΃<���23b=�赊ED����8�v��c�rYm8}��"�0P����b�L��Ѩ�ҍ�L��ǌ�l������X��_t��<�����n{QClWaD��W�] �������x���ng��2�k,}�\q�x�0�h�12n ���/�v0n��9�� ���v��S��;��(EE��Vԟ�I0@����1�ڮ���ٶg���H����:���;�\~`���F�!�6l	eŉ���ʻ^�6�~]<�96y7[b��HE>F#n�P����=Z�D u(�c�oa����zR�����	�s��В���`��,ܜs!��vނq�%_�9v"
�Uh�C!,���꓂�`���r��(�O�϶�1OGz��"����^�9�R~Pp���Ep��#����&��J2v�	�j)�8<mIgd]z�O�Xi2����Egf�;2pOD�'m���)YbJW����炻���'4��5��M?�)���m��lf�!�$
�D�%Ⴏ��ld�E�2k������m�
�E=2E�I�Qp(�$�������*�h:"F��05�� Ye��ͼ���Z�#�/v)���oJ�T�5����Gs�~����gl�����#H5H_m�[��H���_���5��PLP�~�l"p��6�o�::�u1���q�5k5���d>Bq�#ބ~�|�%�^D��O	�Ȗ�r^����̀��k2X��a9y���Cv�~ҢAo?������KF�j5����]��6�e�0�f?��f����/!WK.J#T��Po����x<�\F��Y:6{�f�bau=d�34��r���&��/��^�{'_�s��(�J�7�E:�`��Y������"��lC!���!9QXZf]n	��(��:g�h�������T1W�Ws`B���	�����ؐ��r{�0@=A4��zn=V�Ӎ���w�$uйP �d�x����'���DJ�^�b����O0�/uj�
띄P�;71	��?��~mp�R��������?ߜ[-�������h���Ա��).=�$l}���d��+B<.����?x�
�`�n,`�i�]���Hz�;���+��\@?[����"�,�6⠦�-u��%Ɉ�Ϣ_C��8�O;����3���]���H���%�	y_P�rqd�����!�W���M�7%�W��,E槣z~��)w^�w��� �|�v���[4 
��a����F�D�M}�Q%��R�lP{�r���l��w|pZ;��r�evRŷ�R��Z��]�̤N�(L��ߊA��'ktR�Yd���$����H���nR-���C��1L��^XlxVHYEB    fa00     8e0��p��j���څ�ڊ����?a%>X�8�FsXLS�Ɇ΅�b�u��.�aDoƻ�p�2��S!�g�kK��}�'�O�����3�؝�EKŽj�*��y�ٝ6̯�s|��{)��a�n�L/Ը��\�xg)zo^���%�3� X,�� Q82�Kw���a5�?Ly�:��6f�=�SK�d>�����/�=�� ~e��)�'�y�7٢q�C�I�ّ_e�$I?�s��G�o��[�"1�J�cg{�%Q;z�O����8+NOJ[y��L2��P�E�_vt��,Z���R����	�y>�Jv�L��wV/�]_4C4�l[#�♯��k���g�W�}�<�y������g�PDe����uA�b�y����( ��ed��,��tu�\��a�\���u�a��k,�|�ZV>S��$�ͽ���c_DmzH����L�N&��%R��;��դ�n���P7��O�p��:,�h��ƻ��V�+S[!�3!�S΅�I-i����Dxc�L����Z�'su�a����¼��7A���n�+R.�cQ�(�@^F�+��mXFE�W߯P���C�+�5��>P�D��!�͠(�t�Ngw�$��Pʐ��X�`3av��VA�L/n��'f�N��r��*�4���_�۫R�!����JNO�����i�;�E�f�� Rmv~��c��t�� kC�sl����uˮ/^�j����2��7K�BEV1>�i/�o�,#��,�C�$:,����#�S��3`�VƄ�*�,?3_��^�n�`Y�ޫ��9����	E#��0�@<@�9�
��(�G�{��*��n��%4ǲ���ô�Z�#�Xِw�$}-=П��T��7�f�+�$l�W�`.��\���ʘO��<�e��B�-�@䭏ߥ�i��4'����M�2>ʠ�xaݦ9q��
-b����D�\"UF����u�9�h��/����|TY� �%����:q�4?�B�	%��/<u_�q��Zkx��/�Da���K�+?o��2�\0 
,�d>�C��;��$�h{'��2�a$�������Ad~y���
U��9c�H��#s�D�9w-#*�,��0@&r�P���J0Ʈ95x��D���1�I7�]������C�9��z�J���!�k��P�R#����o1]U�-�=(���S��D+6���R�r������S�������I�3TP�b��F!��;����is������ջ�%�6���$Pik ]�T�����-<E"��.,�Oy��剭��o,#dp�q��nW6�C��"}� )K��>�F�V~g�4wP��s=
����z&lbI���r�ECOg�W�,�ة�.r���A�6�0���Pz6���)gC��Ц_���Z��q���A{��G�ؖ>�L!�_��#PJ�bc��mj6�g1ZoGI��
�I���i��NK�����e.�d��F�j���`cܚ���X�}C�J��3'�6hZ��#��7���� E�����E[0l�.�-�U�r��уx(�Ɔ�m���P���p+���k���uT�Նx7�� �[gPU�\��;��y��OK_����NYY�R��̰�<u[��#'z�i4=����
�f��[V� +�6��l����|1$�_Tx�i��$K}��/hS�wQܪ��Zw�:���W�S��p����	� B�=+�?[�-zCQu�X��<&���x�C���2��d8U^_�V7���SM-�pOȏBR�#戾>	�����;%�
�����L�S��aШ��̲��"v*|��{9R#�O��;cm���~ƺO�%$�E�L���ڜ*o��[j3k���f�, �#��I���o�z	�e]�]��\��`t�˱����-NY�q�hy�G.�T9��+G�(��eP�%�N���������(:&9�}�����=�>�G�0�b�V����&������΋#��#M��Q�����L)�S�*~��+ޫ��.�g�~�T�0���+��ݗP��f�2>\�;M�����:��d�T4�i7qJ���h������ ��;)@�tL�z��9��T= $7)NWu��]�bn��f�d�-�}J���q�T���w1BE�t������C��e������I����b��^G7�����*�j*y��vF��x���\5<|��A�ɤ~�����o��%c�4!=�[����������D�ޱ�R��d��"� ���2XlxVHYEB    8f7d     7c0]�Q��-��>*�Ok
.��O�I��Epp�k~��� ��E�xל�?�HU��?�bЈ�2sdM�F��ȉi�Ű����g�Si�)�'iK2�z�J�3�:�\O��t<�w�p�^K�/߷ �'�6ކ1�ډ0���7�P�W�t�mt�;;���{ ��� ��������Nپ>�Eni��F蔑�c�8P��P�y
Y%���@D��	t&��Q? ��$��'��3�veko����F�(L_�+���z3(�����0��A�sl�u���Sa�E���3�P��UF	C��C^'��2oõ�Su[��-B�l� ���@�7��~r�ʴ���{o�l_���</=H���wDX�=�=��a���;�Q~.�S�m6I��'�pk!T�d:���6���*�� O\�]����,?϶�{kȔ�uk:s�7 �߳ � Vu���&���V3h�Oו.y����ٌE���E�^.kU�9jp�_x���,Ӎ,g��"ȝ�󷴴��#��X+�'���S���Uh����L��' �)m��qޗ����JyG5�j�e����դ&��~��#Y�6ҋ�sUӱ�VL��.��%'�R���u��Ώ�ّy*��
�!BN��S���Eu�=�O����csJk�7��?q�q:&H��*�j��X����MA�]c���,�S1v���/%�֦ �Dx^CB|��z�G)�����S?4�?�rt]o��Yb�x�h��?�a�^�Xc��^��ӻ~��r�(�7��5�8gh�,�l��:��i$uÌ'�����ڀ���]q��-�حZ�KB �QN��4c���ij��h�lq�D�p�}��jp�}��MǱ�tJ���O��~5����꙯[�W��A��.뷞˗qH�����Jx������u�q����	��W��0�`~Μ����banRh�����0&��1Ce���	�gWb�j�O^����}�<��lv����&S����;��b�"U\p��#v��������ƪ��q*!�1}"��u�4S`�
�}�~�K�z}a���O
��p��g}���3�O�~��-��DT�1+	ر1��o̯�G�����mc��h�z�̀#�L��%enL��� 뛐�����[��+�d{�PI��$���c_F�~�7��z(�:�hr���E;E$�K�D8�ɸ	(�,J��#L���$CL�P�Y3:n�|��P��`�\��&c�U�l���.fBi�#�d�ǲ!,~�I�x�;����pZm=6FF��a`�2���}��s
Ҟ+H��<�z��V���~=k/���Gʝ=�LĘx㝓t��>��mXr���31�5U��l��z+��S�,�
5R*�I����3j&녕v�N�F�� ��A2ǩ���0���y�z$�;���^��G^y����J�J�f�Ռ�=Z�Z�R����}���ۿX��]cT|s� |�-)�L]� q�y�)r���b��g��w�ʍhm���8r�䝠G�4Xڦ��r�}��9�n�8Ӧ��%�Ҁ��2j�d�٘p˰7�Z�1�$[�4�+���HYł���g��.ל��T����	�d@".)3D�Ժ�f�`�Gv�1��CT��]���)��m���n*��A���[�����/mt�3�[Y��������hM�	2��cUV���{����iO^U���������N�n�>CtIʢ(�P��z+|W<;�S<���4cKJ�+���FȂ`!��9@Y��� �5�Bl6��0�-D��h;8�H��h�����;�*D#��f~���%��$������w�ls +�2��,������";������_��&��?&�/Ф��Pr+���#\�����x�=g�p����ylv�h���'��$s%�Qw�����������43w��֣�|ja1