XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ݔ3����x��喘�P�&k8ҏM��RO�(�o���M�rPu�[!�I�L-v��N�+�Ј��}HjtM'�PFxIń!�0��H�'���Y�r��D�u���|^?�2r���L!���U�9*��tK-�YL�7����c@a�|�l v�#�j&n�j$��.�r�K�ꛞx\�P5�����O]����2L��JZ ɗ�r}�t+�pUF�f��8n����v?<@�ĥ�,���"�P$z�8萶�q���xr}~4
����J���`RUL�H��צM��]��Н�z��3 Й~�ɍ]�G�8yV��p��ب�K�� ������(�R��ת%��E�w���u^�°bEzJV+|kZ�G�7�D�di��5 ��v���	�]���1���;=�w��)ﳚ��ϖ�i���_�3�i�z�(�����A-�&�u�0�u�X����i�N{?^}��A�ŵZ���*տ��k�'�)�[u�tj��|6�$h]��rY'6mۊ{]m,(�]h��bSҥ3�]EL�H���TC<�*��i�I�{h��0�1��3�XaD-V�8��T�TJV��O���R4�h3*d� U�B�c��Sz�^��|+C����$1͠���W�|+�̑��䣜"X+c�@?�\Ɗg}3S;�S,����t�&�������i���8z�)dӷd�o������s����%O�(��W?�z���N䈅�Yi���,/���+F��u9��XlxVHYEB    362b    10d0N_�W7�Z&�e.�Q�;�ԕ^��0�3�zh���w���f��?��Ր��
�T�Z�"E��T�hr��I��f+c$�&�T�V��<�rV��{�b�ZudN�<���RL��B��	2�.y���:�Z�}� |�������&�M��d�'|�ߖ oۈ�Q��������C�T<��<����	SA\6����j^��Ѧ%U�c)���k3��8���=�>��*�>'��9bo�	�|A���yH������8D�Z�Q'��)�� =bkR�k$�Ɣe��b+c���,��F@h��nNٵ'
��0��N��r��<�}b�\�ϰ���)�����-t�80�!�E[v��.�:ڕ+���'=��!HM0�CDSn��&�q.�I�]�:(b�����#�6�y��e�unqjl}n3�����y��_�E�
�;�����5a1
i���G���t�CxrݗL�������G��?�C#r=��6\n����ly	��L�z�"#L	MDV½���D��F���B�Û��}�[�~a��YS��Qہ���#�xf�����j,b�X:A�g��WE�Àۍ3�A�l+�a��SY��_������E�n���R酺;�#RK�r�w����"�h���BL�~�W�.�T|c�i@m��1����Q솓�"�M^:�ရW0���Fb��M��YF���ZWV�U� �Kkjw�1'�W��x��v���R�c.]���3���U��O�B�vm+R�7��2"�f#���'���{�*�Go�@��̺w�<���6�C�*ė:����<?���Su��U��/%�i�bK�b����n�������6�i��lS���:s0;��i��E�(�m�k�͜lC��>����E����b�@��~���V"�`��:g�Ď�=�n�]v^��:?S{�i�?�F��f�6/��h�8�b�Eu�R6�I�0R�1tgFz�B��ͽ),���o Un��\�b��a����-���)�׃�;,&��z����˷yU%��[�@IAK�\�����Y��C���U,=����"{V2�6����W�}9� ��s15�����	�s|�.S=t�_���e嵉Y$*)�Y4�6�w�v���]�&6�@���p�'��������2e�WG�o�	�SRњp��qd^�3���$�(����Ect��o��{����������խTak9��̬S���׊.l;U�
�QI,V��
O�Ny>:%`㜖���d+9�B�^+�mOe6��Fښ�}��ȧ !Jt,-P�y��
���"]b�J���
��D��͌�������W�ߞ�A1W��c�Us�<�� p�+T����O4�ί��G��ɮ�WHe e<ask�a��Yj<�p���񨑤��{w��8�v'ߋ{���4�ԬN4��sk�<���B�auuE)��݉9� L�/�#hq���O�#ݱ�Nz�����.(�t��)̤]�`����a��e����ۉuXE��#��~�n�Wr�%���z��E��RAt�-&>�n��_�p��9U+����)��|�6v��4K>�&J�.�7g�;����=��5>~tSɛm��!&��F	�ش����a��}?g,V�[T��Pܚv�4��a#O�r��[έ)%��+{�T�� 4�/�F��j��rX׍Lк;�8����%���ev#�	V�����Bթ���X7�Xq���c%}|��L�4{'O��
0Ee��2:�=a�=�?�62� $��`	ć
���3r���9�Q�g��o�2�u<��~I��ά�+B9nd�~��K����V�{I@�Z#:W$1��JlNd���}5$�s��a��\����X�j�2�h�`����%.O1�k��UZK<��TŽ&scy@��b5�3r��(�x�*�t�<D�/0֑�\෩ '�at������9���q�:bTq���̐E%t�4���'���n%�5����"I����H,��Ɗ���Uԗ�Y��Ng��MC��f�od���k������T�E�%���n�f���3)\�����<�J�������bm@VvJ�iܜ�"{��.^@�1S�_W�u��Mx�k�����pW6���0u����D�� ���~�X�ӦW���筒�U3e���T�F���������fP�R��i�;�1��r��3˾鬲���KBV���y{��r������UCpÉBN�pu��ʈ=/�.�nb鎥�6��Tb���+S	0�1"�8����2E�b]�����G��qh��5̥�F���;Ou�Jx��X�[}�=�K��A�E����B�L���i��7(�uͧ~]-����^ ��y��}pME�9���d�{�9���
�Ì�E�I�nC��V�S�U@DD^9�/���\t��/ùSQwt8r���D�b��2	�;[&����������)�h�_�͖v�K������O�p�k�@Ļ�O_x�r�S�u(͈�6N�Q��o�� %���[�n7��a���X����"���/]��2�0�7�:�� B$hi���>����a�1U�D���AP^8� \ډYd�'�ͥ/��.�f�Q���2�* �N��.�1������r"��3-lX����<��#��f׻՛�3�m��R�v����A��	fX��	ʛtR�{C�+x1�G��~R�. � ٻ�	��YDjQϏ�!��򇣨���-Y��t��Ӯ�p�	�����>QmchlԪ
+��ZkP��`Q�-��a5$e���r�Muz�1��`�%_�b&�+5ZA�𺪯��x<�)�e��&����\� �l������m�O�@�r���w%`�,u�y�鈌C��v����K�2�C���@�uNa�ׅ�l�%�hΔoԷXR!�uM�LE7µ�i�s]N��Q�߳zL�*B��慰��JP�3�	�li��S����!'��8P��/�|sV�+���Ŗs���Lz�-��%��p�J��$7f��*�����������إu�D�9��H�͟&����ꔎ��
c��֕؇y��b@~��^U�is*b��Z��e�Y��9��m^q�O��n!a��p��M���>����UJ�	 #
m?p���_�30U����`T�أ#L>�ы]�����t�ʑ��j�:s���i$�!?�T 0�#9?�4��E��2t�B�bvT+�a��?���������#�B������׶Ȏ��
�c}�˿�1��C���ۮ�HN'N��8�����[��)@���&V��C��=�6>Ax7/ƥ�7}a�-~�J2��"�f嗿�2>�G;���/7�����+��'o�8�����C��~�@k�H�c�&�$$ʝ(xGSڎz�Ӆ2�kZ#�i����5��"�52�,M|4N(��&'���58pB&�}>SZ�w�A�t�lL�H�X����	��'��)�N��~�Pz���S)��fRNL���؝	.� ֽ���z���M�:��)��	��-D��������1�4ҺleO�YN
hГ?NY.:����ܫrw�X�r�j­x~Y��ㄪ=�po#��*��+I�5�J�G~ۿ�О��/hk�h��6�lCT�����
E�u�{�Ё����M D��2�������K4��C^�s
�%�J�6��J��Ԋ˥��/!&���I���	S6�"Tf��o���|<�!N��pHN����j%����3���k��!�+耿m�$4� �z��Z|��KZD��U����,�b����N�Y,��.��rb5D�~���t��0?1�/�{��U��э����Pg�N�n�`]p�}�zHI�L��?�o>p���E�����(!��(0 ��E��vQD�֋�mq�LK�)O�~�x�!B��2X@�zQ"�~�Q|O���{;C�}Pz�X��ڀR�gX���pjp�}����b8���7"����F� �a��!}��]�;���K�:R��8ɣiM|$oD�~�P%���S��p*�E�*"��#��E%2���=<T*�|��U	���6o�;\L�˱;}�D����2��]�I��no����%�c�����j��eǢ�4G���Kkz�v��閎�m�5UG����qW��kć�w���^��E�p�7+_��v3��2