XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��W�p�K7Fy��m��\�?��@ڸE.��`il�)sa��v4^b�#t��
�F��7�z�1\m�V�Pb��z��u��n�sz�7��TN�� x�ȍl˘��Qгl*3�l�ŢO'��|��U���O�ͤ����BY��a6�NF,�z:�
�s:��f%�A�Kn�ø~}L33V�Ua,233w��]=_��#ҥ��Ӈ� �,���pu!=�'�~�ı��m^Q��r��R�8���������Sy���-bڎ���P�5PA6�ud͐�48�Q'�]ڑ�h����\X���y����ʐuՏ�]м���x� ��~I�t�f�E��<��#G��g��ʐm��U�'y8�.���d6`Ŧ����Z��& �}�g�|� �[N	�^�)0�\"�t��L�����E���W�c�����h�~���y������s>*~�Zy�£4�����]�'�F�����g�Z�7�Q����t���W��N8m���	���|�6� �4 ��O��?U���[a��-'�^�e��X��\�r�k��ފ�xTV"Ϭ��������i8PhX�?J�@����e&�Dx4S]��$D}����~�mT=`�!}R(d�O�h��T)SkTi��[�a�D�ԖT5��F����83O/�~��fj�u��x�ޱsw.�'"&/i>j2L����5��ΕZ�d�S�[[��2�h��H��%���� u8��;��r�ު�ؚ�!�	�%ۨTK��D^����#�gXlxVHYEB    4a6a    13b0��p���@=�MW�a	��lɘ�>=��8H��n�B�}�ܓ�Vƍ�e�u%���`���х%s�T�)8��9)v��Y���D��涆Š�I�)g���B�?��`���zJ�ߝ�:a��M�:�&��9�Bp#���?3�����r��Ė�����yj�ߘ�A�<%�8�A�v��I��/@n����b1BP�U�5�������� ���u��2���C� 6ߍ�:"li��(��Л	2�����_��0�4� �7���W���d^_b�Z��b�)]y���۰��qV�s����+�S7�/�;W���J.�>v!���En'N���Y��9���䥥u��5�#�0ЫI8������!����YpH7@�$0���5�����K�ۆ�������s�d)�gC)y�� �ನ"ʓ϶��T��3n�,��l=�RK]��^{CrTw�;�͐q��j�)���*��bE5�\�sRm�*4r��G��Ypq!떒�T�t��r\}�GA`��
&�U�ĽF�6�_�<k�:���B6{2���X�|
���[����e�lb�a6�a�W�W�ˇ*�{\m�E�L3���L�r�]�p!�
k6D&��Jy+���$��K1�t�y����$�r\V`y�S��w��+0���b�QB�.�g�zhoXb��W�.����L�;4��x�i� �m�`��3z�Y�WUے�Â)	���]W�A�A�`�;��m��!v�$�\s��/�I(װa�%*2w����(#��{����X�ć6�%���h���.5g,��Y|v���O%����Z"�j��X� ;��j���)�	W�$�W=r��|4 oa�@/�l������@��n�kcjjz��ф@��t�Q��O�O~���R�\b��nY���������6�a�3��~�HO�D��>�Ї��9�i��՜�/K���n��!4T�&�ꐺ�֢E`�Է��mY��{�D�@ͳ�1�㧼'�D�c~.¹�~7�wQ�l��r�[_�<�S5G�e� �s!9�A_��h�.v�|�脎jVO4M�Pn�j?U�(J��x�L��ݛS��Z�u;qKN{�J BBy�d�M9�K������|u���@��E����p�.�$b���.��dޏ؏t�+
}.�=�T�3�9Γ2����ʺ$ ����x�݅�~9����x�E�	���w��D�d�a��ȬX;U���#3�t�!.4sO��V'�\���z����y� ?&%�������~�2�3�/wSv10�4��k	W�V(��e��?R֖�O�f-����+Le8}���s�v�)Z�4O�A?�UÐK����a'��=��#��g�c��f֤�Hjt�����~oP0)(u���WAp>��쒪!4@4�r"+Q)/���:)�N�B?�;��eI)�ܬ�*���)�4/�.iSZ�׬t ��7�-F�F�A��F�ݼ,�#�K|���U�)�	�F����*\���:d�����KZ�(ؑ��_)����1�}���G,��-��Ov�@y�{��㵱9W&�X��?\0=va����4�a��B��Tr�Q�?��<�(�R�^m�W-}D(0�$����m����l�w���%C��,����!sj��D�J�Y�����8�!~c!ɘ�$�uzbԚU	�i3��e�D&HE/78�P@���kݢ��u�$�ȿ�����
�4�r꒷�?��>ʊWwk�=Tx��O�v��gE;�6]}����0r�|S�"��e��=3��2Z�D�T�L�.�/�����sDC��C�/���Ş)�f|�F�0�H��%x��=���*�f�YMݬ��9["�m��9:��_�
����t;�(/�8#���8��%�^\�0Ǚ�e����*���f��k^�%������./[-�2|�ZA]�X���|n�(���d�$�?�yG(A����BO���QB�XQ}8�ܾr�hxCa7`c>���ᒽ����ֵ�)�O�Con�x��dn�W�
� 4���4�W\J� �D�a����DV��e�FX�GI(|v���ǝ�������D|�i�d�	�e$�eOzC�*v�B�7��L�/�;�,n�9q&�o��e42�(@�����rfE����R��:}�iX�9[�;e�[�*�8���+�,�[����#��8N_ރ�)ڹ95�6�>'��(oJL�!���/���ؔ���l�?�����#:�RH�u��Y�H���NY)%�T%GL(��U7��* ���wB�^x�!��M��G�/�.+4O O�8���	�l>�����>s�Q�k%�F߬sE#K��J�&�	RP���AH���rN�~���h"�Z�OSfq�E�+8�,>��T�����c�xI�a]`��б��)�����<X�+�6>
g���5���y���U�Be�q�	�Nh*���R������Tr$�6Ö{�"��I�1V�{K�QL`w󀍰�>6��. �^o��i2�R.��u6���~s�?sG�|��VVy��L�ڀ*����d���@�C���RN@�(�)�7�V�'{a���W�cGo�!�04�c���h� ���=�����3�p�τ�X85��������=z����~�V�a�ݳb;�)	h�أ�8���k��I��v�a�T�1Ȋ�����-7�s����� �O`X�-.I*��r9iv�S�烌h]1c%�a����S�pe(~	2�n��/7	������$wdH�,x�u�����(�e����n�S�BLC�f0:`�\�S+i�^�?�RO�G�]B�7ꆱ3R �V��h�u!Rw��G8�\���(����H+ ����J}�=`��n�(h��?og�0K['�2�ʹyzP��Z�^�g��бcG��j�@R�_�}&�Z{��j�9�T�^rv��a]�D-_���5v� D�6w�#]�t&s��dBA��RG7��Ɋ��F钪���+�.���G�����[�1���:��7W�Y~i�O|�2%D�͈�4����+�_��#l~�7�{�b(�)[S���'��f��>����t�?�Jw |�� �*����D$�l�1��ڧ[M���mx���~H��`fX�U0���2/�:�_v�Il��H|��Ì}���?�a�y�o��m��O#b�*4-�z���s����q��� �yT&wI�3��aǕ�+c����+��º���1��(G�%������M-� ��H���6F
��/�ߊ��5��ܬ
C���S�4�AX��1�!�[��<0o�]�T�h�_�xn��IR�LP���$O������>��N��:���;�c�妠v��l4�tPZR7�"�2�3�Yi-�'�C@�:�G-J]�6�D��V�!��39D&��%�σd�]]���Zҗ:�ʄn)�����g�ȍr�WN���ά�z=��뢶5�hp��.�C��̑�
��I_���+�ɻ��@~�wɓ��4nќ��(3F�����3/�L�s�e�`�����v�΃�U�pN��MV��L�ϐ6�+����
�hh��倈���ѧ��q�v���A�]=K��Y Γ��(0����}���/���S��� �|?q��xw	�0�-ܦA���с�y�bwG��7�!��vd��@K�����.'�H��k�4Sc�_��-���h#G���U��\�����Xiu��jf6�2�j�=f�?�BPQdx���]P�r�s�`�nW9�q��aQ���6t��kQ�������W�h�u�B�pK���e��-�S6����+�W!UBPC���T�	�6O=�1h�Z]�r����3���j���x��Z
���zk�)^st��R�j� z8�ךn�X�Z��m�
�hL���-��Y�{�������W�"I]�L�_ФR���L4?q�Q�#�T����7��r���E4�GCۖ���nF�_�$>���&/���0��,�!��)�']�5��6|-����'�e�-a��Kr�Vr�4б�kľN�����2,>Κ��q1�����v�L����;���*5O�(�@H�,�}U������i^�H�f폮L����kW�Tջ��Z.:ڻ�6xHD��'{��/�B��4���n�����K��I_zV���������~K�{�O�%��z����+�M-�y`��w�Kި�>#י��b:���C��ߔ��1R�@5��B��Ɗѫ��X��cZmњ�S��Գ���X��lnx��z;�GW�S��
�&�*Z�ܷ�� �6d�Q�� U��q��,��Y�k�5��eu�C���3�T/�	�}؋̸nq+���ԙ?�  �QɜK�/3CF+=�$*��/e��T�+�_�ś���Պ � @*s����ɨÛH�3��ڢ6�֣T<�埧��]�P]q
�ܻB!.	����܋B��b�d0 �Lg[�6�Z��k��Wgo�Q���v��E�tG\+C���d���8����<!3�9�؂�6ԏ�»)�M��0���n�ؔ��a�鳇���5j��Y&�L�	��c�!z�ѫ R�zÓ|T(�t#u0G��UǮ��?r�௞�}�W�����bR��pzg�af��>>[�������C8�_n�|ErKL"d�_�L埐�Q��,G�G�����?;��-.�6md$�N!�]��?L{�X V5N�Cz�@����Z�-W��a�?�v �QHұJK����ye����şyj��cL}oH�D[�x�SNܩF��)����x5����>��ib?�P��MA�l����6�b�7���$��W����9�7�h�s�'���C�<�FйB�ݚ����Ψ��)!QL7�/;f�kk�,~\� EQ�*T�Ck@�T�K������Y��j�i�6r�ᮚB��>:��*�����ay��W�