XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���+c@�����o���抲:��949�:b�z,���m�����s&��;`$����έ������р�SIrW�\�3x��ޝ@�yI`�u{�
�Xa@E9����Ӓ���&P�7\5��߽�v��7��K^ir
�ꔦt�h�2� ��1��J|�G���L��@[�~���r�P��kk6a�U��GN��+J�����:.ƥڹ���r�b>+ IV���h���~%`���y�eH1{����SX�g��E��}�K��������}бwɅBp���ƴW���<���q���Ni���9y� ��1#���K�)K̦�b��6O�LD_����7�iV����Ϊ�<рq{U�x���b��@.��uH�G�I�F���O(�(�Ģ�᪆�A2�q��T��ů�[�Ir\�;%�t-RS74A'�u��
)c�n^�@,�"�:��c�0l��N�,�G-|���T-��0�+E�~�Ȧ�{�ԉ�Q�0k^+��6)��)�HDp�n6���I2M�O�C"�8]+�u�64�!9ލ�c4�����yN)^���S��������z��\�x���%�����P;<�]S��3/Kt#<��\Mq��F��4����dM
8EEn��L7�t�oA����:_2�����'k���߸v�ۆa�T[�1�k�$�-L����Y�r�(����i��UVkp(����h�����������嘲,xA}��j72�r8>�Γ
)_�d�09�A��c�h����XlxVHYEB    7d76    11a0ų��O��[ղ��z3B>�j��V�I ��2l΂��,�S�D�EUТ��f�R�z�*��¼�-����7A^H�޻.I���������aJ?cND䈅�J;0Z*��#�\�D�N���U���v�%k�m?�b>��{׉x�;�,t�t+��4?"��胨wEtA��!J5P{�V�0�{յ��PGo�cLY,���ʖq�ˌ��{{�bI
�����ޏR.���c��6�oT�/����6N���3k"��$4�R{R�^-&��9az�ۤ%��l���Oh�2u|_�tK	6��9�������kPr8��}?��l0������"����F;�_��oЬ��G>�D��5�=�?�y��ܞ��.�-&M�-���}5.L�B���#�QD�A���c�N[�^7�>Ȩ�[ˏ�_y����}�nyG1@/��1��\�ws�,:M��`��`�V���_C�OBX$
�8����]E���jV��n���ʮ��n�$��۟E�h�&�X+���u���4n����X[-/���0t�#��mViĴڽ :��ֱFX^�5�TC��LH���	�6�N�]���dm���8%�R��<k�:<��j9���ތ�U=�E�%2��I}��x�)r��֡_D���8y� ц�Z�����TQ��. u%��Ȕ��p�jL�F@��V�6�'< H������\��">qb��[<n��$��R�>U�bQ����XH3ֱ�@��e��AK,��ߋ"_�^��0�?q�ٞi���B4A�6��d���^�T[��Ow�.�p=Ve�$N�f�ւaIA�2[����$[W��u�\J �2���_G}p��5�D�!KR��y u'�>�����F99��q}����"�*'����2m�EAX;$���JK}�^�,�\~�6%[uO}���s�-]��w�����A������α�0a!�4E����]��{Z�5��`COK��r_�#W`�r�B��*��>k�ț����L5�}믦�iu���Um���$S`3��8A�{�i���t�lT��39g�`V��'7ۇ.��\k�|)��(Q�V �*I�xh�m�<9��uǮM5�ki����)≯����f�W�^�Y�p�\��^��Y�X��g
�tє�J�����S�~�^�6�fw��u���=i^�ծ�U�Z���`<��,�C_�������B�*�*����������C,�c`{��zꩠ����r?�E�B"8L>(���'4���h�,�υ~�Q�]/�d�yt'��������W(���4O14E?#8���|Ǉ˰)w�w�������.���@W%ͣG�Ɣ���ט�#q���k"�8q'n�{���ܔ�ʴ��{5�V�p�K�ӆ�S�m�0O ��Ə�����g�*�VO�r,ѶϹ��@9R+�%R`�d����E"��z�n�ZC{������݂���E���g�v�e0ߗ+��.L����uLe�m��̾��Î���'�t�Jx�� �'5����<��+��~�X��f�aB�A�Z��E�+�K���}�)Qp8�Wk˵���s��3o�1� w��j)U�g�����}��5��r����'ō�;
cB�d[V�F�Jp����d��ܘ/���U�/s�s0ҧ�R��67�P�?���3x��~�paY�/��8 �:�B�h�Ȧ��Qa���Z�,�X,�_=7��t@��W:����ݑ�C�R�Wp��\y6ߩ�'��]')��.�Z�6�p���n5�K�2x�׃q"����u��������)��cj��p]�l(��{�﯍)V�R�Y�k-��<9]���oh�d;�w��3��e���!?Av�|d|��1�m��_��ѥ��m�x	������ *q�j|J��n&��׳d�W39�P�Ue3����G׍�|�\;�?��u��)A�6ud;�4�%:��o�T�4�
�M{�e��mA�%��)*C� ��<�������$`�G��6��l�9�Ҕd��3B�4{�&��GAJz�0��Q9�ua0G�W����\�k󚮷�����A�$�F�!G���t��l�A��zb�Dɉ��5B�(�ڊ�nh�ּ�%?��Ff}����AS��"*K-��DE��Jgg����|�J���]�x�zZ���/�P�$eqSV���U�,#N�t%��cQ\�af��AX�5/���Ґ�~��T.���X��������/s�АyTId�v�=6�⓶��"�4G`�ɩ>���NF�
��YK>�F?Q ]F���7��q9�'������<�5��N�5(OjT��*2��`��G� Y5*\))XH�60v�p�UT���W�v_��1V�����A_��e.��$��� X�[��OEˣ���*L�8�KgG����'�9����K��q(Sh�J#�8b}ۦ�r8���a��E�wuLȔ���6���ݵU�ѿ�]��)g�Lj�`���Y#��N�L�x{u�\ӻO�G��t���w<(~�b3&�=�9: ʀ��#ߨ�8�c�/b�?p�ݶ��z��	��*�ה[>(z�g:����L}n!6a՚�_��d��%����ƪZq�×�Sf�n�jw���k�S�m��v�����(Դ]��Ev�+U6cD�_)vz�6X7c��M�o�r��R��a$$jp�wr���B�{s�'p�M����ȂY�WX��_��.'3��Qz&�~5���*�|�o��ks����w�b�#�D+�D�K�Z�ڬg�Y� &Ӻ���ͻ
����o߀��� ?�H���J��c���
���yR����c����W��}���\�s}�`�C9�a��~��2�Z\�4�|5b)*V:�Ο�SKX���W���?���B���qBGku���[#~�*��C��?Hʄl�R�xtp�eD�쑌s�k�7�`��;��{}�(��5с':ƈh(�����ll�(��Ş¾��!�75�7��<�(J�EⰜ�8�g;��/���^�n�)��i�9�WB@<�M ?���&�vv�}E͢��/�h!@1�Fp���k�]<&��D�8�;n���� ǖ�D`�Tp.ѕ��@Z��p�8 7[�;[��=���5���?a�>��.�Ot/�k�$I;I6�s�� ���z����M$y�.v�!�\"|j��j�ų��!܌���h��W��֨�͎:RP*![�Y�M��>���	I�B��O�6Lv˪<�ƌG�'��K+[r=����aX��W��a�P�����5��h*n��3Rm�nŚ�@��!=��f"*S�B�I���ț�7���A�F��Y��� J�	��GT��l
:��#cr��z1Q�n��f��Χd��@^��Iu���:'��z�g�>f�r��N8
}��	D{�fSe9�ߓ�Z;-W<q��K���K�:lJ�|O�9����������^z8y:{-�1{u��Ar�`�����WM7N����ȆВDҚ�[��Ŷ���#�FN%�ӂ��5jbn��*\ԇ8�6��!z��
5���޾����i|�3Ӽ�O��m�'s
+Iȸ9�U4f!�ۚ6�d���z�U�k��!49�MR�಺���f����p��y(�`��ȇ6�7ͯ>�̮&6|̈́��&s�dM:�F��a�ݟ��T���B��H�)"] �
8�{��4J" 6��lC
t^����$�p >={�3H��Y���F,C쌊���;T����"��䑥�������)_4,iJ�b�L��.��b)w�VE�-+j�VBG�η��Rݤ�|.& &x�F�~xz�e�!_�(#mj,�½����ţ��7��o�M�	)w�X�{gC�G5n�K�\|����Ο[l��O6��NXP�,�&���.3:�v^����d8�"�^C��I��^ÎtK���ewE����T�w�Jw ����E���l�a+�������N�[�u��?QYD��V��T]Yeu��(���-�#� ��[� 	�h��o,K�&ތ�0��TTvƒG�I)h�U�	z��^d!���L,H�߬�G/��jiC� 4z�^ѯ-������<`�������תv�!9�]Ļ�7rQ_��-�q�&������"��/��.E"�=��֔�ۚ�
�"�t@a&���:���� ���%��"�)��ɪr��D/I�i=�R����J�*��1�A��QgL�4�kj]�W��g-P���C{I~��kjaG�g��6��{A<O��ț�E<j�����%f���+,Z�y�Yb�s<��V-��D��$�Ѿ҅RߋΧU�J�F��mC��Ó���\����:�J!�~al��c�Llޟ����Ai��֦Ž�"��t}P2�V@�P�1	�Ke������rD