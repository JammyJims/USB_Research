XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ֽ6u6W���繟��"���c
-�m�qn�.����� �߃�&!�:�)�S�|��0K�`��\���"�Ń�mXA}��.� �|L�8;x���Imޢ�é�}!D�E���A:�C�|^��$!�-�8�:^l^���A3�uCz��e8��o��o�,�J�;m���KO^����a��п�R��t�@ޤ6��d=Lϋ�,��f�м����	�Q�hE\Mf8#bp�ƵA���$���d��l�t��������5ɯ*�2W\2�@^�D�u~���H_h�ƫ2�.�y�&uyq�������}�ԇ�e�d4t�K��3]?��9��!)�Q�"-�����c�{a[�i�!/�qت�Aw��t[3��&�$c�-��q��?�?����4`��fß��(S[�"Ws{�!�br1D���^��?cUɚ��}F�{^���4v��h�,�5V��h/~���X�2#��z?2��터�V<ed��H�jwv�6�\\�Ϸ-��*3#0?]N���n��u�r�N��k�g�(e���Ey�c'>�p�7>���Ǻt;�tw���{�����B��9ϔU�:0k�h�cA�1S5�-�.K�+����H�����x��U5��B�E��)�1�yk���uw�|��i`�(í����Ю�}���R$}2�m������c��fO]��Er\%|��+I˶��1������}�D�����H+��o�Q��*l*�[�&�o����y� ��'�O!�����XlxVHYEB    3912     ca0�ޗ':�>y��C�4K�\_h��� ^�y���}���2���9(��P!�~.D�ܣڥiI���r��ջލ�`#�6s[�0�T�f ^Y9˚��3��lŝ��]f�X�^i�5p�@�S����Wр	r��/n1�����z������U(y���'4q�љ�ޜ�t��1蓉�c���,�DAu]�ZjC9-)/�oZrw�~jS0�!_8v����=���r�z�c��,@Z������1���6�9	�{��?��_�b��������Wnk
��ěgb��ܤ<���*w1�/M��[�~��S��.E�a�5�	����i�F#�#��t�O˗�ufH��j����f��<9���[`%��릷�Z&>��i��c�&��AB/7,�M1w�#���M--�w-�A��T�J��^g-d�ݴm�n���])R}�GR;1�Z��-�t�dq���0�!S]�deNou�����b|�wLln��_(4��z�t�/�Nω8���M����*D�jH�&JǊr���R�&�h��~K�<�F$&Q�!#��#O�.��P�\S0<������q�j:�y�5�<�-��Q����>�e��a��� ��fL,��.j��HҔd,�3u����>�8,��D ��N.|��Ɨ����ۦ=X���1V�0���}4��P�C�jF�Ή��T^:*�?���j
��SY�/UVҶEo����Tژ-J�����lUE��j����
WG�($�Qf.�s�[�Μ\Q��O���r�k�������ykȧm�����*C�`���t*��L��,-w/;:�`#]Z͚zَ�Z�Wz��̢�r�%PB��:If��ho1�<N�#����q%�d8~�X�d��\.[��&�![,&@����<��d� �g|}�+�w��C(_5���Q�]�G��6Jdw�2�۟�l^[��H<U<���j� * ����,�N���	k��-#�&	(��\q�,�Qb� /`����R3�������G�>K��EǛɭ"p��r-EEu�NR�l<���r��k�]�8�HD�����6��N{;���fZw�ۼ�\�x!Bn�@�kp� ��8�����6)i��<��<��㾨U�{�Zal[k�F���L��{�n�:T�Y��nf�!]�w�������r���.�߱�C��nUsd�>:���6 �����w���r宅��xM ���&HR�T�X��zހ	f�~����/�Z��WY�x�N<��D�&B���-Dt�u�	60ϴ-�!��P��L�H�T�E�R@���sEt`=f.��@��=ò���.Y\���C�"��җ[�CY3R�@��z>kl1����9�8�թ/7&�w�����)�R�!1C5q�H����/kI��~l���F+N�ڸ^�������p��o���4�Eʊ��1�_�q��ks�4�EK�Gi�|y��;�����IɋŃ�gk���i�K�Ę�C2�v�.u��_�$<ё�ul$FJ�GZDr!1�BW��U�v^(����_�Ӣ~�NA!��)X����\��nc���Z7��z���(���0a��r:kڍP�}�ģ���
"���y$RﷅJ�F���|�Zy�^���D]���W��k9�Lj��f/(�T,hǭǠ�U������^K|-a��%Jf��I�j.����ZK�ؼ3�����ȁ���jt��s�K~�k�@�l����C�E�O.r�sb�!�x<�Yc���.	�r��.�;�W��~���-�jH��KA�OT:�������5)�e�65T�p�s�H>(؀�����*}��O�\�b�y��͏wt�|�>���KO��GV'.�(�Rr�G<��$�*�.�O�Յ�Eş:�����I��F7[�l䠟h>t)��L���rZ���ŷ�d��m���v��.N�>�O��j���Na�ÖX���k+�Z���Λ��-��Q����/��I0������O�w�K�4���9��Kk*�(e��v>P�
�QL���(U~[{��#lNg��s�z?ޮ�b.x�#E*�a�9���E�1�A ���G�[��F-j���]J R�� �^)���\2��2.�,}��l�S�_*�� ����:�2�'1F��H3Dt�NR3���ʊ��E���ӱZ��!L�)��Uke��TZK��oѼƼ=�Z��FheQ^�&1hb%G��j���K?�Q�w�g�Fde��ey�l�u0M����>����[?C��hI��k�#`{�&�6��+W��	��u�}���\'k����}$$�����yܚ̹�8)���3<< �nF��#���cr��=�I[��$^0te�����Ҥ�2��ʠ��`[�^.��É�5V�ڒ�Q�r)/r'̏ ��J+���Rr�c�_{�b{�әU:S,Ϭ�iӲ��(�"�Q�pJXjƇi�A���W������kۊ��R����CA���`j`{��3()6ƌ�og��r�Uv����B�[�@��=Y�A� >bW�1��tUY	0�Z'��~ݟ���Ȏͼ�ԣ"Í���Hվ	�����ox��(�G��Ʀ�A�Z���^�r׳i��ŰL���^#+��*�LD_�����ӓPj�T�%��;�Ǌ�nC0���Ĵ+,�bH�Ԡ������Ұ� �:鸶e���Qlv7A�r�I�M��Ÿ��>��ܲQS.�'�e���';c�_N3�'��Q���0r8��	n�ʻ�U�_����E��$��H<�ȶ=?o/Ő�$���e`hO��<������#{4��Y1�|y�M��w��l)��<�7�Fa�ۖM�8��XR.���d����I��I��K5Ԁ��E�A�ٓJ�R��&ڼs\I�a{�1�np��w}o4�V8��H��F�� �����?��C�\��]�}����LВ� �A�E%�����d!?�:A���敭Wͷ��k,debwq��k6�[&_��e:Q��ɼ4ȱ�a�C�̚�5i�@,`�3F��i�ǡ���L��C+D��V]R�������5��G���y�'�b8�^c?/W��-�.%�tc��u����B��U��k�jVVj[��}��W�*��ޟ ����u`�����j|��/�P�`w|�6!y�Vb>��2���u'cY3����8��5���z4lm�