XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q���u~+,�p����5�7}��r(�g�EE+�K�q<�f��B|LD��]���C��d�k�P_ڕ�N�<'�º��v�Xg�\+A-���@�����R�/~&H0!�e�4]w�B�B��y����۟��dH�5��z���y�0qz�Q,�����N��
N���c��F$����"q;�n� ����g�ZI�O3�Q��#�BY���|
�?L<dT�It�sFŨ�X6��(Q�p�SzC�T����Xv�&P��L�' �G�dX1Ћ��W�[�����:�k���	l�2� �Jn��`7�}� ��`;MgA�Y��+�1P�N�����綆[�t݌�y�/�m�Z��bA�AG����w/������Uuq �S�}��Ҷ�b�[/���>��3H�`�}gC=YSI�`�8�3q��j�v�PS����j.B¦���r�d�0@�s��0�61J7"�ƞ�k��!M7�fyڛ]0�v�VoC�i�J�9��X(��(]�Y�f?;dJj�57�(��\�ƕ.EտTE�U3�+�q`*|��O��h�L�Iw��u�:�ߺ1���TdH=Y��VYaY�%Z���=�-�����|m�Z��j��W㏫�2!r�ѐ|���)J� +�e��Zf�_!!w�ϴh�~-��y��e>(�a�*������W�Ђ؉�F�F~[I���A�v�;�j��O�n�UV��>+�7+��U�lȊ`��'��,��[VӐk	ī���yR���kjOCH���]n�XlxVHYEB    fa00    2970U}ƍ#'��y;����:\��i��O�#ͷBJ��^�����Nu8����*#������H�Ί�[�Pw� D�[RP�*�}�$D�p��tb�QM�]�kx�"��z���Zd�EŠ�C:�����R �I�A�uX��Th<F����7���M�R��2z�k�_��M�0˽�]���8vdwZ:�L!s�{8mKR.J𞆧	�3{�	��f�:�XD���L���.�H�]��g��M_bD|F��{#Z�4�a���ѻ?B��~"X��*d�&�& �M;�y`$�\~��/��si��KO	!�Mk�D|k>����`�J��_���)*��p����G� ����U���C�{�*�l�,-)�ϢO&i��	��|�319l ��Ӯ8M�t���b��G?����}�w���68!<���L6.x�^r`(|OY=�[����:����/�Ei���{��H<V�j�B�k�����&C�I��PV�k�]��1�rL&�gg�f��O�b�S@'u�3�f�U�I�c>2a6��0�i���4v��.@<�uN�=8k�+�5�Y|9М�����9��쬐��OWwNQ�M	)\�����>�P�5���zF��'aCna�:��#�w��L�-�Ȁ�­�"(�t|�6�~��£�<�.~V$��$N8�&�i�����w��]�a�a1 �:[ �n
������?Y��U�I-1���2�~6a�n��mY�%}X(J~%xc\xk$�ߗi0	��g�C|n�n�\A��Q�'�T�����C5�|�g�n�ʍ�H��/E_\P;�Z{;��]%�Vt������Rk��lN��p�m��@�����E)j��%�|dK��pV{�M�����b̓ج���S'�ƔR�51���������=|uԐrGTܤ�NΡ��o���λ��У���7�Ǥ�3u:*����Z�~�ڒ�+;��Y%��&��J�
�v�3�KʯG��ݕ�G��cg�ks�Mr���6���2a�6�8��}�@���1�m���׋��ܫªi(0�P#f�8�m�y]S�p�6,�ږ��_���!:�q2��'�|Ay�w~svB3�D�$9q�̟�,ˣ�=Gǧ�� ��sѪ�����6%��؝1�Y��']�7����0\����w�V��'��+�%%�c�-�fe�yQK�ZԽ�g~��K�[�j,D��!g�f��X�_كU��;��t�Go(��Rk3�
q2h�f GoM8�L?0������j3��=?������z]"1�E����U;�-��DߋA��ky^=]+��{�i޺��1VLD��y0?A���-�a�x��3FW�b�.������/�����Vl��b..+q�|*�*n�A^��TF��˨=���U��@i��V�l�<x"�"-Fq3L����.��$6�UEF6��m�V����V6br��P0�q0���YT:t�S�ߜLW�
z
 �V�re@:�� W]�⼌��w�1}��Mc��濞�~/�Iه/��4Q���|����H;)֙��Y�w.��[A�&����n���$B�J!�!]��(���K*2�]�w���>`�U)~%���Oу��F�����i�������C��0�N�¨���${}�s�vƏ��j�@�(	;�����9sN�;�gmx�+x���s��l��g�RoWL܈���I�?�r9se���U����g��X����~8M�ed�ԅ v�|��r���t��y7����?��6K|H�Td��m�д�"=��K�]���S��*���S����5�T	�w���������u�+.SC\�%g=��$���ʪ�bcE�~?�p�AUڒ~��[V*��T�$^{��*h�G���;FK��On��iU��她���Z�E�ԮѠ��R� ��ys��ꑷ{m��L���q������ۏ}�7pX[+Y��F��}�����7j��^yv�/�U`l{Il.�^џȂN����}�q�y	M�?˷�$C�0X��^��ͫ�Г7/�K߬���u���n�kb���,`��v1ϒQ����m.}�)䝍`���� �)�34��1�]���J��-�����u�K���hD�X5����i�@��C�9����rEE���]6��w�{ r��wq�(�S����~5u�d�C2_׼��	*�*bÉ(�>$:�z<z��0�6�~�P>o���
���W6�"�y���7eۖ�ǈN��'��(4v�Ж�u��TM[�~Q�M��;�X���-+�]�#�����[��D��F�1޹��a26����WЉ��a���O��b(㥖s����* TK6���}PU �͠��&�A�x�A��m�㣖���_��!rC����N�R�o ��І�@/\gO�<��Z?=2q��[_�\��*>qu����9�)�ԮA*�N!����������0�`QH�(i���@��[�/�:�ૂ;QZ�2����ݨ��%a��Q�[(Q���l��3\
S���a���1��۾�A�V'�Σ���Q��HEN�`74RV@�t�}�O���ŎZaO`u]jJ��l���[pN�0�s=:Aw8ۜ��i�o;n�&�$g��\i��Mv0�Ůi�B�Q�s�bτ��~#y�d���
7�Pe←�\���l��ũ@���@�����9 %j�0���s��*��_ ���=ᐁ�.���᱆��3�$(���f?�S�ŐU7��q��;2 ��jC@\d�CV��w��/g���z٬�RJQG�P�_�q$�Trg��WVC�*jNwŃ9���n^z��1��L�+F�!E��Le2�ġ�);����)�?�ع��!���+��Qwӆ|�
E[�ø.�	�pnwc�D�����,���*wÙjE��� D=]��N7���#m9�غg�bqR��E dh|.5�� ���Vyd Tq�d���]�]8��\A[�w��6R��v�^K1�5MV����*�[���	��"__�u����K��pE3j� 4�_7 u�@ڎ� ���<��~NU]�]�C�{`U����3��"O���K'��mf R�c���1�e믤����ww��O���������t��?3WiB�^���Ϭ$�Z�늹���$9���wBo�z����k�&2��̉f�Ô'��9_��C�Ob?�׃�Z+�-̐B~UCƉ�����!� th.�u79r�2|��*A�f ��"��݀,R��Ý�o-iżH������I{�/I0鼁A羶�7�n�os��4��ϳ�R���$�F|��)F��Z����h0�:r� ��U��y=r���\r���+��#i_�88y��m����鯠O��X��l|�6o��a�G�#�>�6��\�̈́�Et�f�l�'7�p��V�S��������%ʧ.b�1'�I���F��7��Ia0f��L�3��<����]wN8��@ϿW�Kc  ��6��oKZ9H3���Ա����Us\z'=Pq_���!0�����g@��e!��Z�����[��ϣ��hn��0��	R��qJf�.���X��}�[z�)�[H��C��n��Le�ט
:
��p9K5�nZ��+#Ec�����=*��+���ND{��{뼩�rK�U9����	����2���,R�(٢@��g��k�l�����-x��3��E�p"��T/4`ElS�I�X��=�^�T. ���{��bDg4~�:���Z�$�s�&�.G�1��4��
z�!�{(;R��c,S��5������l}��G9�ڜ2[���l52��_�R�n�~���ȿC���z���0��D����!��}�>�UZ��>N�I�E��ɳ	�����׵�2 �H�N5�M\ƚ)�\}��I6Nw[�"!BQ�H�l������p��@�۞�6Ș�ZIo!M�A��X�.z�e$�dǡ��'�_-M�,Ϡ�K�q��5���4������r1�H��s[�Hp[I>z����I�ym������<6l�TS:af���#�!�[�
�		���!ͦ�u�%�o�_hs$�9!?�Ö��V@�}�zj�{�
 Q��^�1�����F���H��0י,=��ҩ�����h�-!@^~W�Κ^���t���2�Raһt
��K�ʝ�P�/Z�Ԩv�@�����@�QWX�ﱈI�W��<�W���d�$�Fb/V3r���3e�ӡv�Q{��@iv����Q���S�g(q��#�"����~��c^&9�}�ل!8�ɕ=]�f$�X�+0�[Ey�K����u]�Xd��s8���ڼ�sy[k��6P�E�ҡ���!S��(�h�;�G�YgUz�ɛ�:��z���n:G�.R��U�[;���^;��j�*`�̠�������49��@ŝ�����0 �,K�`��Ć7����C	J�˕8�������G+g��ldn2���nŜK�9P��WӼ��	��L��Q��G#W	��?�RL����������7-p�0�����}��遼)�ٽe��0$�9�*[���7bYj��M��{��b�ݬ�C���[�b�y��W��?G����*
�{�`:Կ�p+������|��q�����-�I�6�N�3��Z��m��� G�\�3� 6W�=M�����pC@y���'֝21��-��%T�� ������:��Y�1vSKQ�B�;� ��Y�/w�(��x^��8k��y�yK펑;�P�}�����U���t��]�$7�G���.�g��]t��g��� �{(��i�Q&?!R~U�v1~'b�u��u.ǎ9z�,TM"_ �8
�����_^'�Jm{��gGgưD���J��Y�q}�E�\xD�����mv�,=��n��6�&(��\�d`�n���\:��{@JL��S+B��f��f��E�"˽��������]���pj�֭u�6-�KP�t
�ȩ$<�����ܦ�8� Y��|xy��/I�*�+Y�!�U��3M�xEqZ�p����r�:h��Ń���u�6��0@vU���c~_l*���u|��;�Ɗ�7D�0f~�m"�Y�#� ���}!e`���&��!?j�H���o�]s��a�a]̆1U� ���J�*Fҽ�%������IN�H�tr�ĕ;e��ݶTAVB�7�p�Y��WA q1]��:�;��	`�Lϡ���f�4��vzi������-�u���������O� ��k$L�a�����(�jŜ?�&�-y���I�M ���o���\�0\��0Nd�����_gl�M�Q54.C�U*�O���(n<��}����f�������r������t�n���%0�[Df����Ac��y$��G��SPu��7�O��9uf�ږ�D��w�E����|�~{'��b�W�����V��XC�¾E��BG"�����a>iZ[�����V>�+U�_�^�\�~�F5�~���OO�"J4�@�;&B�PP� ���Kw�~GW��O�����E�Y�ؾ���3ӑ⋨�~��K�-��Jr]c�����·���Okbܙ/F���X���8E�STwh8dk��;1«�Bn�pi��|=� �Wc��?;��J��e����9�Q䏦�f���r❔nk��!JN��'���c<%)6�y��6I7���d�s�
%���y��;�Z���u�~�~xtM��C�N�S�S�5%��]%���6��~�l..�b��*��I뇴A7Bf+�?E@�C�����P��O]�!�#�݅J��5X}��!G�iU��r@Y�1�9�sɃB�b�(�)|�	�,ȩ�HIy�=G�t��������>��鍶W����q�g�y��"�s�z�N�~�T�@:Xp,]�f��ʪ�V¾��6������ꨏuNd�}�YU����#��	�	��FU�i�}�'�I>���_���F4�0-	j�'���Z�Y�D[\+��Z#�(��� ����|�rM�*A���V�e.p�$�:�|i�_ͼ~�h�8k��p��h1��>Q�Ȇ�YRu� TEc�?���=
����,��\�W�H6.c���+O�����p����An�mS��p/���R��d6vR�bj��hcV���[�Q1���?��R�פUr��y��iR������f:���{{U(�������h;�d�*�ow����BNa�����ÚF�S�6���T�,��o���؆��ïx�~��xT��e�
��� ���(Y%KRgT���.��2���W$�5��J����!���y��p]�6�p��іX��^2�u�i!#�f�x�3R<ԥ�6��ܥ���@+Y�b�����f�����eYu�+�B���@1��[¨O�pi����/��-�m��s��D,!.oo��\c(5��XaVhU+�bVg�Y�A�����[!�He�x���~��K��X��)@��$'I����W���GT����U�V[�v��'wЉq1~ Ї���?���?��,��FOS�u��V�L��Q0D��O��W���T�� ���&�_���a����1>�a\���t��d�B�s	F���I�}�5���3�iy�+h�;����B���c�������'4�z�܏'�L�
Ȗʰ-�,�)��3��`U���A��_���|�J�D͡;�;����˘�y�*�l͈>�i��
�*"���e:��P���
r8�捉=�[OSZ+���)�W�E����)s� �l��Z�"xɡۃJ׌&[�ЙBK�9�Ɨ{^5����7��6M׿:����%�y+�ּ���I(1��_ݺ����H� 08��C7?z��1�v��9��+��y8y�����lA
��zl$���(�aNP,OS��L���lL�FG$Cz��q����Mʙ��8R��we�y
HkF���ڬ������gݔA�H��z�{�����U3�6ߋyP��V��c�3�q��o"A��h)J%��h&�Aj��Qy].���D���\}��`��-��=%��"!�_�;��#��o]L?������	������6B�,���8vd4{(�p���!�(w֝4-=᭼Z��Y0Ao�[	
���Y$[O�櫏<=O��΀�D)�iC���op��>����=K]T�|�¶��J�$>H����֝��%V��iǡ稕�FTхŪX��o���y#6���⾌���e��_f����5ёW���(�G{�G8����Vs��4�'��g��;z�0
�f�L����rm��\]�L_�%�|�|��n�¸:Rc���P��"���ptZD &Y�G�� �������a��� $ND&�U_46�[×�`I����op�c?������+�F@��7c�8�*�Y~L�D2֡h��4O��9�5m����g}�XB�Eɦ���	�GU_��J�������W�hOtsZ��}-,��)�yW�3)?�^��R���~�$t^�ns�r�hc*y��X5M^��/�}�� ����,�IH�����S�^hv�6?�������N��>�,���Hs}
L��6<� 7���f�a����lE}��g&G79��a�hY��\ӽ�
 ���T?d�G���2uR�L����@��\�+Xtsj��7���z�ȏ�v��(p��bXѪF�Fh
D�jt�K���^�������#��6��0��)�oڍ��޸�LcO�7j�n�� ^/��:o�g:�q3��mgaL��-v̂H�-`�> 7)ٕ�*���{�Ry�3
�J��vwԱb��v&c���(�$�/����[�,��۹�,瘌�w�=9�+Ox^��-N{D�����?m1~��F�J����H�|^�'�O��L^:,&ص4��~�6-/\Ou�,���U8��-Zk=�l��9���f!5]Cq@LT��O���4K�����Jle����/@�"[w�iн�(�I�Tw�Nچ�]g�`ȳ��!?�A�#���b"S��;�	�Ŷ��)Ëw��~	p��'z�����|��d��4vZe.af�q2`��Ǒ�_쿍/��[`uiE�H��Na�2 �p��]X�Dܜ:+���,���)�=��`�:3���)��l��R-x�B^��?�� ѯ,(��(�'�5�K�oY
0M��|�Ro�?�c�>����*�q�R�D�N��%�)�3#�d*(�h�B�ɍ���Vv�r�ࡅ�76����fM?=ͷN7����F*9:MTvʅ�N�I��c�:����N�M{17ͨ���7����#�Yq0����0�&��nr��`�A�9D[����j�ݸ�Bށ�:㒽0F+�ol�*}��T���W�~�4�e8��Cd=�$�C�����������w�h��UT���n4� �M� ��r\;�H������ёU�.I��wn�9�H�_���r�z_@�k4�"D�b-|aC�N��}��_S���	�h�J��x������o��ԫt��Խ��;y��Ϭ<��$��5U�XV�4�V�B5����WIf�X#>
�����R���&ݯl�@@�_�VX��NYّ�Dg�߈�o��9i��h��d9k��ia*���j��CA����^ouD!��'�j�p��r}v�
)�eͻe�m�B�,�q���D��Y�75�7���9?cd�ဝ�zCR�Uj�0�z�*�I;Ð����Q��Xi`��P�`J�����)��6q�����݋�$�e��F���.���7gyA����d�#p�C��"��9D��G�hR�1x���췮�11F0U�roJ�R����8#N6@�������iT�vQW�������U�^p�
��e��;qvr��/c~7ЌOt�m6��*�ڀS�*��q^�G]֯>�tH�:��͔���%�#�$�����Z��E# L��� 1m�Ͽ; �AI�&�`ƣ"K	@U`�p`�d�.#k���L�d���s�T
�=��͇!MS�S�Cҍ|��Q�
��,&��H�-'��&l0r\�`�C����ԧ5��]&��wLC�c��D�̼�T5��p��P��&��]�p�P�$��b���O�����eH-�I��W6�Ѧ�Z�&����V���u�Pr��i9�qm�����|
ʴ\��ԡ��R�D���k��ͧ��،�3���V��<M�#�M�9�$�	c��z���&^���HYd�D���d�^��J������r�I��R�a��.��3�M�><�FL�wppon�Tw)NA��_���j�2b[=��됯�5��ڋ ���\/�ә��X�<;��ى���x�[h.��0 ���=9ُ�4�3���2귀qd�ߑG>�ٌ��b����â�f1Fł��hPV3�M�0��O�[hɣ�]���J5I��UV����,Z/���\m�蔐*C�����Ѫٸ@ӿ�)'������6�ٕ%�^>E��\��у]��J��j;P� �;��L�Kh�?h�`	�"�ߦd]�!提u�!��IU��i<���V�'K���0$_[�P`-��x<J����*��>熍����=G�n0R,	ʁ5�E��K��Cw�JniS��o������my4��l̑Z��D���ܑ�Uj�;�r�q��/��hf ��uC�.0���p�4�"���4ӄ(�ו��{����ڢn�ثӵѻ0�#=�~?��SN�=�e�Uca�����9(IeI�t�i�R46��	A0�� �:�[N"3�>�5*gL eῚ�����1(�p�0�C�t�j������o;����:�1�u9$�T6;�]dw�ipң�@oo��]gڄxU�&Q�F%ܻ!���$�|�?k|��|�a�S� z).<fH�c.@��#� &����S8k��xˈ.Cl���9ނ'y����DG�؀�5�0���W�B���0|'*N�m�É�P���}>7x�ջL�kKfS����X�^�֒x��|3 �eBv��Y��ӥ���vV�P��՘; q���*���=ߖn���u����v��$�4b5י�7y縿�r�E��r�V�w�� ���q�|�aI ��� �|x�ħB��W��4_-����F	>�z���h��V�'e��.��Q{��&�@��+��^a�7K	tw�ҝ��н��`��&L�@�f���[5;ouC�qZ�p~Cy�Y�Ӂ[Y5�Z��џIH)=�H+��<�e8h�DH����	3��U�gfd� 1�Ec�g 1�Bk.{��L���\5](_�=�dl)�C-�;���$-גg��`�^�C,��[X�NP
J�� ۷�fW����F�}t㽴:Ww`�*�+�&��)��I�&k����>�IՖ��\�eQu�����@c�~xH4,cp䲧���qXlxVHYEB    35d5     a60�<O�.�|h���sz�(�[��^,xgS�� U�8;��I	����f�X I���w�m��:!�n��ψ�����*`zW�DU*�/��-����m�7�r8>�Π��.
�we@`�\���	����ܗYmU!�g<�^�R�$�����
��znQ�S G�,A�P�{R�X(6q��g�\`Ћ)�w�����D_л��؀�\�I�֖V=�r\͵[��V[�QQ �K7�.����p�)8^��o^G�1���m�f�M���~Y�`/x*�&���o�˓�/	���l�|m���1���1�7��Ć&����v!��0�^�M-(���;���p���O-��M����k:�r���j'7f
�"2�����/�i����cR���� �$x}�ʮvѣ��"Y�9}bDCp����o�&T3��W`6/�D��#�B�@C�ũT���L��븮\�w�h�a)�+�ⴤPvH�P�{d���<k�xR�q��[n�
Ɣ~+�j��q���Y�u�'������"�m��'�"��֣?ɏ[��gӪ�bS�sz�(�O'Kj	Ż/�ZhJ���e���n��|^�n9��ԝ�j	���I�h�co��:�>w����~\b^�������5�47n{�G�r�'m�`۴8g�Bכ��N�h��	��'B]��D��[Q�'� ˠƤ7F8��,(ZͷR�����Q4��D
�=�+�x�������\IK:�n[ٌ�N���}�������""������TO�!R����M�QQ���4���'~:�����X2K������s���M+�Ƣ���wv���n�����׋9��N�@�~���|�(bSͩ�9��'ݸ4���n���k���� ���Ǉ�A����140w��b~~q�ݤz�_��υ���7z��k.\�8	1w��h�T��z�-{58�LCf�|���<�<�gT�@���w��W7��=D8w�;��=�Np��-���բ2ᾑ�YY	p�zۭ�4�aaР�2*0��z�t�_|)JZ���zQM�<�<c�ߥT��Fe��b9IB1���mBwӿ`~������M�Ӯ
�T���Ⱦ�ǳ�c|/�
�&SL{�j�����߻����V����Mc�ٶJ���a̴�m����zɗ��1��F�z����K��w����d,�*���:�8�A�BO������'`��M��N�2����٥�.�:��\�jƅ��U�KT���䎜��E�+8�@,�紦bW�2�鞢i��U�h���Kå�fd�)6����C1��Ѷ%7�2�Ջ��l�N��#�ujB2
)����B+�ɜ� �(�=|�O�Nh�4&S��a��tƐ3��[����:ڰ���1
<:&ZY��F8�N�j���zz�X��8����j����yD:���,K8������E��?�nLA����C�)��rU�ΕVh��\ T~���<�J5�^�,m���)p���ش���"�uG�5���hw��,�[3��>��)^֝TÇM}R.-������K�iM8��
p�۹{�\�w��͑�O��􁷨Z[%}-�C�=��,�hy7�E��<�����XL�^P+8���3T��\�aaR�Xk�Ct�N?[�N��)� VU���a�]�2;O���O��X��غ(��(ug!ҁF�˷�U�̸P��%!��/��6�Td��\����r�yt�<�q�Wʃ��%#���
��pA��]QC|�h�[��*�~�JK+
mչk��� g���{k%�xD�x��C��3�Z�K�Q�xW l<����n�!�fԏ��V�7�KS���|�	��k_���|�B
��=́⛝�T7��qR�C5/��5Q���Zq@���t7�6�Uɐ̅�/uM�-Cz�Z�O���A�y	�8��
*n��;��U�n�-9p��c�-'�(��v3k>0���Y�vg��p�ǐIр���z6���C�W?V�Zgt�>&l� �=Ȭ� Q@�gLy%7G�^�kũ�H��ԗ�	�4�#P�������7S���?4����p�:BŦc=X.-���Pa�'��-����Q�0��e�i�D�bO�5�d&�����=���ْ�`f�;��|p��0H���j)��R�u|9q+ߑ����t�����F���~`��C4ݰ?�,����$t��9�F���-����(55�L��E~�/�Rq�)׉���C���B�k�f���l�'��94L�Bl���U���k����~���i�z�m�-��Lٍʨcp@%lU��y�^x����"���S�\�ǝ#�M>qT {]�N%3Q�����NM�$0V�=c���T.�ڱ������j�z%�O"���5`���q�Y�<�L�>�.
�"p��h����c�ղ��,:6c�A�i��b�.W:0|>Ű�h�_�����" 7�Z"����������JqP����9g��������sn	�4}m����N:T!�ŵ�H�����y]�V�Uh>��=M=W������p�����-OZm<�[`���:��Q�+�mfx�G�n�cӖ�xGP�,�H���=,��1���NQ�g��LU�-��u��}����o