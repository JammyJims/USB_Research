XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
�B�g���[��ܯ	��4�8 {�2x�J'����o���խa�w�L���ȯ�]�D�q��; ��"0�A�I<[h�u|g�Y�8�\w(��u�ȌP.���#�?X�B.eZ��x��s�b�f���_	Tn:	|6�""y`���l:�Q�#!�	��/i%i(l"��=.����m
�p���G����0����K(�� ��������]��r����,/���q䃃�H;�?fA��)~�0:�~0���OP���<9j���^m�����qG����nv�����mu��Rܽq���[ V,����oK~��ֈhʛ;�<�#�Y����h#[+q��� X��ԓ���P�L�ir��2Gzt�S�5��,u��ۀ>uv� �n��xp*�`�zyMU����H���F@f7G��@�����x��'�-�LwBN�F���}����/��$S�$<9F�|�w���\�o�'��GH���j�8놱a���|�7��
�\�GϽ�O�p���&ٽe��Q�ԑ�G����̶y��J@ORPՀ�_�.�0������$v�0�M%���zW��<JC3�QϓPUĀ��6���\��_�����A볘��z�+z	�����7�G�7-QLdnȪO)��aD��z���j
���$������`�>>�^J�ZjZ�����R�4�p���N�o-]F�|LH4������og3�9��D�7�I���������O�������1�zd纻3����0"�?|XlxVHYEB    204e     930�-Xe�f�0;��.������*�������Y�4��^<'�*VM`Z��;t�=���qDf2������/���t�(�ϡ/�r������(Y:İ����ʧ���m^����r��'�E��G8!�=-`WQ��]�Ѻ	�"m�9�+q|������?PCd
M�G5\��[}T���K��Dy|���� v���k4��J��<�/`��wt�����:_�1:����gq�v�u8����P%�Fc1qG'��g��خ��?k�?����+]~l\c��3v�[DO�+')U�u6r5�:�,���i��v���Η��5�����=�擾�0`q;"��\�۽�^dt��t�Ɲ�9��-����M�]Z�6���O����ow�j�����G��Tf�JkJZ�;6���EۣBޣd�3��C�ub�=?� ��r�
��-����:~��_�9�Vb�&w�����e?�^r |6�jW%�6���j�sD!��c�;�[/*H�Q�X�i��e��0�9�J�h�@[�1\�Q.�30F�u�c˿CN��?'�k����ɖA9�:���B�MV?�	�Y��m ���Qx�	�c�!SF�6Dc?6ƥ!)��m�/�c;�0����Ӆ�^�ػ�w����k7;��)�����!��"��?������Ի��>`�?o�R	ʉ���G�6�B)��*o����浪Q
�#�j��:����&�n�Q1qÌ铎�E��l�D��M�h������iܽĞö߮TkN��O��|��H����~��n-�L?�F�o��t�$��5���y71�c�5`����=�p�? �G���������	��ь��ș�3��˹
�.}��z/d�s���gi?�Zo� &6��\�Cg9��t!/��p�C��!�8���]H{U�n��AL% T&ق�ʠl�̏m��ѷ*��[��H�2�^��@6
��'��J�Ñ^6m��z+����`�B�MD:t�_, \�>L�C��O�v�<��f��r��q��^2̏ʪ�I�G��}[�C�o��F��zAk����D��α�T�u�j�v�5�Vn4�:�5�-(�[��3���L�R��)i��m��Nρ��.'1�ڨ��e��R����˰N�4�l�qbF� �0����v�щ��̗��(gԐN�qڕ���?��#��z��l1X�Q]���8��z�:\dL���������[��x/��$c�n��1���0�=��$c��\\�y���H�����R�F�A��u���*�}�ڙM������Y�uo»<�������fX螹F9ͭ]Cw1����nc�lRɕ�0_ǭ�#��'�e�%����ټ�2/�h���Tv��B��Rb��`_N1�"�����}-�}F�����#����P���`�ؖ����s0a{��Ӧ��Y:lT(UCW�v�ĆJ�N��ϐV����q�t��*	�~�f�g4Yz+�l�b�	�$d�X"
�c�3B0��=��;x��f6�z�7�X�9P"�V<m(s�_�G��������I&�+4�p^Շ[JV!!A��)��D�<5��ѦڔOӏrl±(��<��i�Tھt����w��ϳ�^j�DX%��"�Z-HX+����y��.�!k{ݠ����	�ђ���l�1�|����"[ٷ���Ƞ�^�o��kޙC���ϙ�Jܼ��2%�����͋w���x�N�a�\�y�i�$�c����*��d�96��B����v��w�t���ᵵ��N�,?�5�T~Q���a��A����/xi�vn�a�y^G��'ˈ�nC���г�����m���{N�_�i?�X�y_�(��Kq0���qL�|���I�) I�����j�#|�w�GD#a�jݑUP�-;��Q���2p�H9qu���̉j���H}���R#��+܊=�ݎ���'0�����$�_���C�U��.�f"��n?�5�͆����@���.�^���'�h��e��n/�� #�z4YG��U��o[���ILK#�m'���묁�0��g���xM�녒���e��5�����Y�	M0o�K�Vl�)2B����~qV
��ڕ�*Ca�=hdY�N�+��
R#�r+�N���qa�N�'��r���K��&c�"9n�������6�Ҙ�CBv#Z��=UKt����"&�Џ��J���sש!�g�ewJP���s�bUR�3&�NW���!�*����Z��b���s}:B��W�}�|�7s<U��i��2�Z���$I�>j�堲