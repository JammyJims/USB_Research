XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`�=J;�#�i���A�$߮�>��]�DP���J�k����~��Ͻ?�^��GY-��`I#�XID.<q�(T�Uz;7!w����	�T�	~Y*�K�2��-3���A���c>�����;CpCH�XW�:T�!�D��c}����MP�d�)E-����Ahh��V��{/�!�����&}��X/�s�ȝ���Y�o�,2ഠ� �BL��C?+c�\�w�K7�i*4g�M���Lƕ�.{���u�bB��:��%�����V���^�X�I�|/z�!T��8Tձɠ�l=���t%�_5`��b�'@&:*\�qz�_���_'(���C;{ٕ����#�����Y��	�3�)��[p/�M�h�`���Z�_�q�Ԗ�Zʡ�Rݘ��?�݂���	m{�Pr�/�(2�q��*��4G��?�@Ja�w���B�,?
]jȪ'����b��2ԫ��Ⱥ�����o�R�7��u�R�����qu�1��P�A���W��'씩�/����1Ͻ?�����$Z4Jd!��ʩ3,բ�\�TY����|�r��#Lb�^]�dB��P����M+Sj�7��s>t�Y�t==z{$T�`�2#̼�Ƹ�O�gف@6��"��Nh���#wg�eX��ވt��At��[ysnq��/���+*����:������^�ci��t��	-�(����B��&��|-a>���sXw��T��7jx�E��&���Wi!�I�z �XlxVHYEB    18b0     820a���+�8���Ҿ�˪akP���P���0KCN�|�n����z�J�ې�a�u�
`��:������y8�ˬ
�}o��>
`L��A�J'ǾD>�|m�#	*�9(��8�t�+d[_YH]�n]���J]l]w�N=��&4xRu���]�畕:���&ԠB�]���?��G��v!�D�J���#$t�rZ�+]ӹ��U�+*���! q0�%�.��
$܌۬��v~n�{A&H1��w3H��i����em=����Pm���
U@����H�A�.���n�&X%�t�)�f�U��4%�Y��R�769yC��K�����>4�����C�*�˺��]-H���b����z%v9FX'�j)����^$�禟�
�|Q�� �x⾩EG]L������/Z���;5kϰ�[5�WJ���%A7�z����Aΐ3Nܻ���Ei��X���_)24b�dX��9��8B2�>�K��ۋ؀u�8�{mq�S܄,�
$is�2Se/��Ԕ�d@yB���IF�g��rrv�����A�V��ʶ�0�4��žts9�=6�D��n�\��n�@��׻a[�Il��G�ݲd��5_��Kd?)���5�����/H]�<A�\���j?��#y��rO��ꠀf�;J���K�=��闐�,̺q�����0���6C�O��z�ZJ���ƈ�
Q��� �U$��49�����$��	��}
�t�S�Lw���v� %,$���HUUA�U��쓁jTD Jyt�Kg�y=U }5�n�W	��ټ�<�x¶V��C��fد�&�^1�0` hd�+<{�1z�m��Q�Y��rp�%��`����)��o��N F�)�%�Íal�=^�uJg��T����� �B\���j�/�	11�澠���oZm��s{�ٺ��V�]�h`����\�f�!���Po������Y,�����WZ@��`���_��F�D! i�<�Y�C�N�B���������4ݶ��[#�D;k���KV�c�,��O�N�����I|����;�6�D�T�Z`�\r< ���u'�`141C�5w��|noG��Yp~�ub���Ճ@��u2���G1ik���t0�y��?S	��,I���p+����ç�%�\�E����9�S���@��W�M�XM�E4�}ZIݷ�k?��_�>�t�N��;P�Yee{�z�d􎊅�ժ���|:G�`��}]O�I��Vtv�{"���cE�o���"�Ǌ��F�a��ݢ3~�M!t��0��m6�˴���ⅷ���KĜ+�F�Hߋ`���� {���ȧ��b{&�_����@5�G"�>(V���ٺ(�p/4�n��B����6�K���w��R�õ��q�6���_Ֆ�j]�	�PANώ�a�Rv�ಃ[���3\ BKHB��~z��M���Ihv�Bi9t��  0F�<��6����?68���]W�ơv�@���F�������W����^'�/�2�j�3��C�5�S <5%#��{���[f�d�$�'��HaLX�p�'�G��P�!��}ԣ-�]F!@)��J�lN��}+��?t4���;�u����\;����Z�]&F��gN����d
��E�}��֯,\�
��Y�Ep�9$����/�%~ɫ6Q��bL��������_`4������ĝ�H��s��Nq?M��8Q����@���A�y��x�+��cA�����%̚�O���Vj��U&������(b���(o)H�$?�Mx�/��P�[���] fv��ᤑ�'B�;�8�?�J=v����Q�5�&�k�"[�n��6�����_'�2�g^5nL	c7�Ph�IT�/�p�(Pl�RAX����\B���y�J�$��o���+W�����\�=��q̾YV�`�	��<7k��>^���[�rf�05i>5i��@lH2+���]4a'����v�m����D�7��&���9?��
k�uVN̜+���$u��+�G��IS�p