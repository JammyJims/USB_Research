XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<L
4��/������¢>�
m���0����B�U��eڕ��m��c��AOB��ޭ��Z�ۮ�������5���} �^��?g_y�>H���gB���m�	>@��}��o'%�B��J�?����]p��"��q��_�k��?_��QWv�Ĕٰ�-w�-������$ ��'�Ʈ��;hg��e������k����g>������m��9�L��k�/ї2�A���[����M\�
�f��}/'���YDA���=1�\8T"s 
Q�f�	�N��8���Q"u[JM�-�6�b�bK�IfU�����G3G�m5��N���_��!�i��߯N�$��0)����'�~_��r8p����-����8�
	�͗
&�|ހ��-�:�BvbS*aZ�{]�͎.WcX*E�G��N�B_]�)u�V�����蟕 �aV� 	�od,kIM�F��7��w񩳦�he��h�T��� ��dV)�F��F� ���� ��9 ��t�R76�.�<U1��D׋̬���:�ml�.'��p#�O��Kmn=;�r ��5G$l�\i�_����~���G��G(�}!�����K��`�{J�*LQ�o�Og�k�v�:���Y_�z�]�}�����ӆ|��]8���] �}k���Q�6K�xi'1�-4P�sI`jy�|��Q|T��91w�d���Eq�(-�����-���)h3iS+q�&rs�ח҇�|��-kdZ�N�Őu�J��i}���XlxVHYEB    3bc6    1230v�l� s��;�:��u�qv� ��}���SH9.`����@��4lw�:;g�ۜ�XU�7��":ֿ+f��W0����t�iO��+}Η%C�
�xd��M�/$���	s��,���6�:`|������ΐ3-���'ǎbya�=l*r�LT��>�Q�9)7ql8�~`q	`q0h����2������q.��J���g�"�D/�Z^�mfI��v�/��ؿ�5�gǏ�����׎2�.��΋�478I��Nj[n1� *��MnҍZ�M�E.�~����"��Ԣ�Q��9�2c5b a h�
m�������rT�}/bp�ت�2���[��
p�����k�!���[�$���̟�����;��k�2}���9�h����h�,��xO�)���c�ʨ���� �-^���5��}��FV�<���5ZŸ��B�h�OV���̀/�rg����Uh�#�0�s�Wh����90���69� �pu�qs��$L�#w�иQ�Ġ�q��9�Х){r�x#�܊y'6�Q� 꽓�G	�8���RE���%4���h�AAIu�1��"d=6`������;�X���λ�#�,6`(/�I+8������6lγX�uj���7�@j�۪�������`��ʠQ����oe�8#J|���֫'��aMs*���c�!��[@$��S)��?�$��c%;�i��{M����^�Cǝy,�s��6������?�U��0����q@J�0�N����څ���&Q�=����]��<��ǚGj{$��U�ͽb ������a����ST�������1��s&S��
�����0�F����_���^�tT��G:����gl�<�?�����Ux�l�C��P���#0z�z�A`+�`'7�joQ��\��`C�E�m��5��=� )`©��(h�h�s�P�8|V��"?0g�����b��U}Ҟ��*���y�^�".��}l�\��밽�A!�&�G��z3��yϫu�0�P���{�X������6��m~�h$�;791���s�8 :S0���l���B&"�A�;mf������Ao�/��|���v��R���
;�ŔClZ��vKS��"̛6WS���G��2G��������pG�����r
���"�Tdr�F��A5������n ��|������]�-����dCfU�	��xU��E}XO�j��wJ��@Q�yJ�ݭK�����Z5�� %7�¿O�4Ve{YAg�Ԫ���I�]��W}_��c����bڪHa�O����:�:��Ao��>52s�����NVx�G�)Y�����6F��sX`#�w��H�$Fz�K�/$B
Q׾2�9����HU�ٞK���G0���K+,8�v�R?7�������J�m+e�m$��)]���ɲ�����:��7��[=��<5��RN��I�D�#��<=J�S�惍�K�e�3D�S���7eIk(b�#�fT�J��)ts�����e�/�^��3z�,s���!Į�a�˶�;��^0����l���
��F?'M.=}\3����Cs�@[�Nhx�\�{��
��e=��M'��,)c�g[���gp��Q���V��{��zF��)���C3~	�I��E2��f ��2��&�|еVunk�ǘ��	'�'�Įß���BUHI<]�"�>�oR�_�����l���*�y��1ߞ05`�^υ������cz��`��5�nO��?;y��%������D3�<�qV)�Ɲ���5���G�o��7������
C��ꨫ�/hq�Ջ�$P�+F�������`��euD���d8K��Ō�~RS��&�_��ORʞYr�bw?Jq���z:���Vx���[�ؽ�k<.���"��|��4��{��x�l���/��ś򜩑�	dJ(��������l��M��F��A.�l��i�yUp���G����)��x����6_�v�i�3/t�}��h�y}8�8(�*�|�6�A+�LTx�19�dy(�&Nr���m�*�i�u�Q��XB�G}��ѥ�[ϩJ,��Y���vZ��#]����'!O�@@)����_D���W�7)R0w��P�E]z�c�߫���qK���z��ˡ�q%�d�l�兎F򷞧(H��8b���,�|9����1H$���D��[��eB�0�ι1Z���q�J������餒W&{r��B�Gt._��7�iG�Ճ�7l����[��2�'"N=�:���.�>f1u��Z��l�E��sŠ^����(�9(v�$��i�#�z�`�O����1?�Y���� �ᗴ�r�D_>�ֆ�oA���>���/��	�迄��Q��M7!ь~�=B����$�>g���@�ְ��u.��w���9߅�q�Z��-����"��V�͔9�~��e+�àf�+%^s�՛Ǉ@x��l��A����@3�9�;�uI|���j�D���s#>�*���8>龾��J��=�����?���x�.��0�v@�CΔ�ξꔀ!�	�LU�C�Lr�����LjO)��!<I��J�gb��ŭ���A��7��8Eg���j�d�z(�C$�X�
/�u��n�ąp�ʯ�(l���3���_�^�7��˘Yb����L��Io4�gw1����;]h� )������;��8S�v6$�T�(�����1�<�TR������	�И�(Չv����P��}�(�����u��Z$��u�}5����C<.��8/.��5�,AU��s�c7�AD3Y���[�y3�;nO�1	0)���݉�S���`j-A;�;%-;~m��#�K{=�G~�m�u�D��\O$�l������#T��=uE�~hK�R�r�Gu�'��<���՞��Q?�6Ԛ��~��h�3���/vɉk(�v��Ї�@}�H�m�g�lttp�4L���\]��J#֍�Al5���5i*�	�dV�P�|ɏfPiE>�\���}Oz�3�;s![[�J_jT���wY.���/�^���u����9����Α������(��=�qi]sS=��(��,̓3��+��F����S���� �kn"PDA�Q����Q2��38o��0gb3�':��i@��۸�чL����}�C|@y&�w�I>�j���./�攧-� ����L�2T�D��CE�c��.� -n��!�� ��-bpPB|�� �=J�n�S<9q����c���y�{�Z��Y��
�BM��2ݬ���\��dɆs� |��4�K��b��\��}o����ʫ� c�Un�x��..�f��!���m��"���h ��@a!Tb(Y��a�-����i��g�X`��k�u� �I�L�9�
 @�B)�!��4��x����*!x�^ϑ^�/�Z�7�i�$���,��~��x���k}K�>�&Q�e�˾%�5wl������"1�࿖8q��6�gՉ!+{A� �[ri��3��x�����k�v?� !��{�߳��`���{�j�����^���I)��sn���jx����+ǔ�s�����}7�����l9����K�t�D��H��#fqg
kj�oJα�
���u��e`��`�y�L�m�،+��ex��kRs���7�ڷ�:�ϻ�IF�оK���|��������YX�R* ��X��s(.�H������1��%�����X����DQS��᎞�q�䡒��w9*a�L�buk1
�Q�^T�@E0���Z#S3��ar��ѷ�"N
����Fe`0��ǌ�����Df��6�:�ST���~�c� O��L�=�9.X����@l�xJ<`�׆V�΂��Ǎ��@|t��K��;�d����Qٯ�gSv�ow*��4��J���p'��,s�߬�͠�;38oMӎ�_�9y����*�1�\�t���Hw(�(˘O.죏�"w�2H)��������3�1�D��B�ZUib��D��{��FR6뱑�qh�
$V`7�D�[�yWI}O���V/���2��o�����ݧ�ԷSaٟ���H��Z&Q���X^��/��ƲP P�F9P�_UqǴr|�ᮺW
@�r�4��* N�ք�a�h�W"���Gt�V�ۼ*�_�qӠ�������w�Z0;���JV�Vk�*±�*��"��xO; ��a��o�z꽑�k����=ttq)�Ӕ)x���^nV���u|�%h����U�zC_L�eZ?i.��Ԛ�����?���@w#�35<�.f�
+��I}F�W�e��m3�q�[T�ɥ�(���Js�=�
k�F��7z�˖�N����f/2W��K�N����\��'��jx,�D���� ����]�Ґ���r�9!���p6�E&����R!@�JB�)B�zE���	�6> >T�+ȘX�bc�BU�@#�u�-�$9�u?Ξ�L踝����tBU�Q�,�]䏘�J�R��b1(T�����!x�K�P`�l�F�Ô?�B�%�F�N	��tV�fT�R�ik�h�B�����Eݮp��8=6��J��D�]ԫ�T��