XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����k8��=��6���k�^��f���)' �yR�����o���r� �z>�M�8���GmJ�D���V� =���hC�8z��B��r3V�;	�xR���J}�^�@��M#���+����`�������"϶��*����a���{%fp���[7V^%I�lf[r[����	S��K8\�HD����u����
��G�/���6����x��;G�^��J�[�,���~�R8��?OnDu�s�F� ���������H�p�[�����3�>�F����2\>�-�Q�S4�
|�[ğ�#����B��K'����"�N�0�
�ߺ�t]���72�X��[M'��WX@|��$��v�-=5����M��C5�?�F�C�v�|��`o�u��x2i��7ma.�ڱ#n �PE��܅v�VG�@/5 ���-&�K�������O6��؝�v�(�x���J���7�6c)�3d�6��$=��`O򺢪2(����S���L�͸/�]��(VN�_�<o�a^#��]�[ԾX<�\�x�(~�S����9��5m����M�
'��浉?+z��&h����SX܇A���o$kt���2`�`{mFd	?�s�QΘg#~�WV�V��<6?{�i�_s? �g@�p�0�K��y���3�i��7�eO�pe
��u�톯oI9���ϋ�Ÿ01�E�ذl�KFY�x�1�U�M�G�� B��c��$j���,.�gqe���+b�=;cL������(܄���XlxVHYEB    4d24    1040-o�J� >��w״#��������[����q����i�ĪNޏyO�����Z�y
�B������������ꡊ��d�YQ��M^;�p�_�4fh��. :�A�f�����̆���ٕ��þ�n��[�&]1��Ï�<8��x�YKkv����ͨo��q4<��9%����A��\����X�(��>���p���6�V��.1����Q�n����E*��}�b�" � r�PeF���ok�*�w*�g��W�x�HN��K�]�����(7�����>&�j�*��aA��ӌ���	C��(�&n���/����v��!����7�+J�
�l��˨`<���=��h���ת��=f�O���F�k��U^k��?'j'���G=B2�e˓+%ѯq�{�����`-қ),F�HRr*v���@4(c���}2�F�jZ1�q_���u1��l�!jB�0r�.<~~����̏�����~)�R�T�^X����(j]7{� IB�:>�9�E212R�NRP�b��a��}����܉��x�hl�Ϧ�/��a^�]�}���O9w��z!vT�GZ��D|祝�#� �fXZT��#�n��҅I�R6
���(��@�63^��maN�0����@����ty�OU�D4�[t?^*�d5))� G��� �ܑ�K\��v��4�p�����C�売�S��;�0���>��-��O��0��!\[*-���ziV��f�B����Ҭ��ϤQ��P�h�Ò���o��qkv5JL[��L?�OjiP�8Q>&2L���ۿT��m��=�/������F�*�\�Z\���k�[[(xG���Y�-���u̟gT
�I��ئdK]^��~�djNN�zx�iWRSIf�0	���y��$\(����a&}/��K��b
��:��[0�U�-K���G3��>�r��n�.��HF��	׌«P���]�CiW�[/���w|��k�բ��AO�r�����T��Jf��^Tp�X����n8��˘]�l$��d�G>`Y��Q�7Q�jSN�N܅#��5�I�x/�5T;���I ���y�Z��Da#�6���x�u?�T:;J))�Ѭ>�\%N��������):9 ��)��&,҇
>3)�A��*��)���_慤?�2ǎS��-������Ň�j�Ϫ�Ƹ��"���	2-�o"��X����FS��?-�����=�\	4����*k��sm��3�v���F�Յw���*�����+,��,񛟱����� Br߲Ln� 	�(01�{*��|'#+�σ�=@,��<t��;�Beg��a*�~�X�Ζ�u���N�/�����ZŻn�h�����%�E�'���'Ȅ�)B_]gSM��i�Ǉ�i�>!7����0T�5k��k�.����&K�F�EQʤ}�q�;�PW¶zv��u3�Q�H��=�NV�f>�Ŭ4s٠}�
�7���=�m����
���4ys�8�)sGZ*�Pg���5.�P��\Bii�nv�֓�sx��1CTI�骖��d�
��/K�day'a�gM�_�g�js7��J�+��\�ȫШ2D�Z��E�y�};[=\C�4���-(�����|J��F�^�6z�	��m�����G�/�MXT���6'�p�x�fcر��͸x;�2u�G�p�
E����7���ȁ���M���+y�T(���͵�Uπ��_M?�M紬�e9E?���,Jv���:J���:?1�rF�4a�^?m	2�\�`�bon�f��o���5/Oe�a�}@�u �������km���eK =�b��ɒ�F+>d?���J�1y��K��|L��9��^�\�K�!����#�ΐt�:�%Y�0�XJlZ��}DEۨ�tw��L���Y.|s3���=݋�zz��anN_m�pYŐ����q���&��":z�_�$�!s7,��b:���8C;y=���|ۧ9�@-,��/S��V��v#E�g�u���\��ؗ<&?2`+1!�m�t�H�N=t�HZd�= j�=�e�����DԺ�����`B\�=�_�L*����op;|Vк7!�dV]��F�}�5Ӹ�O��6���euV˩Om�1�0T/C�:"In��c��x�_��K7}��]�X�\ߴ���
�՛fa@rf�O�/���?*��?/�U���
A�r�m�0���b���Ȧ/#��~t�H3�]�`��'��.#ux±���Hmq�E��Јtl[f�U�Ȼf*@o�D�0Y�2����O�"�;$����huR�G�K")��:��9=vx�T��w�ἔ-��2*sUޫ0O)&Ė�h!yaN�=N���bi~��Q�A�����eZ�!�V$ȯi�LI���o]��/�h��L�t��c r`�H�X�횙r���x���Nb������UF�$���s�r��/n����xF�tjaUs���^�\�>��ɝP�F܋抓o�&=�Qߤ�v��l,�a-����$9xO?=OYiֈL�SK��K=xn�k�q�5������� =.Z{�3����@h\��>��x�?!��o-�ԛ�?��z4)S�#Dd�y,k? _�[Nӫ�
h��v%��48�<W:\�?Y]4��?�?�)O�Ʈ���W'�ٴ�b�p9rO�KS҄yI��K5����ɗ�I[I �O�C�Т�W�E�g
o�t��	*�f����$�����9U7����8��W8�/'o�p�U���y���1����jn��p&}����m�۝B!���S>I��mJ+�CO~/m��$HB�(��y���~^b"��f�fZ�D�f�k۫��������uKA�W�*� ��݀�:%EJNZ��2w���V�i�����aL��ݘ`-I��Ce��^A6a�C�_/�2��b�|�i�  Gf���t�ϕ�7���d2_��t8
a�/��ҽK�,R���8��D�M3Q�j�`�a:��n��b�e�����8����-����]�D
�Q)�^��a,��yh�H�&[E�����[S�?wW�^�2<d�d(li:$���!c(wio��{`� x]
k��J1�����{�s�q>��ʛ�9��5"�����,d�?D���}C���|TY$ڥ��Gb�Q({����2�J���G}���h��nz�v��koUn�vF�ƭQML��O�R/����-�����K����j��_î(� `�[�Ͻ��{@>9e�+�u����+N?���iF��%)��b�R�3��2tZRys��%=w�p�D�o��ߺ�)�v��A-"r�`Uen*}= �Ԧb'����Q��u�W%��p���w�6�b��7!��]��h��x��n���:u<Kj���yw��k𣮡@2��R�[x�&�n�Q�+�8	��s���!E�6�qу8;�Û�c��� 3k�qJ�|��"��?\���ڟq��m��=l��58ޅ�*�/ͪ)SRѰ'%�W�����R�*�?���y��t�����Vy�3CSM��;��Z97��*|u3q4��c�����Dm�*�%B���rPI�� ��)�t͞-��O�9_w�؈�Z
���oR����[����y���T
9{l4e�a�z��w�����ۻd=�Xs&��hP����M��� c�o�o,lG�e�Ts�'��׍[I.�|*d9��RA}�5�	#5�D���O��f�cu����=�i=0L� wT�ZK�:Oj)m�*��.P�vu�/Y<Ru?�R\��~M��^�`�(��|��'�8å}�j��e�i�iq����Օ���9:�^,i�C��Z�{+m�4>6/�bp��Y��l�J�VuAT{\�����_�F��xe>+����]b���+�䉩A~���^}F��EEyI%E��Q\�Gd��=����·�$g�Y3�ߎv�fߢ��FaPUtx��c��f���9�|�Ws}�4��WPB0PP֤�
.���i���D�8��`.f��PE�ZJ�Dw���c@���<ҋ�>/B|7j����KD�|���\m�)! �)��7�	ܠ�2�P�=� _	