XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~�=���Y%��Y�/�B
 ",3x%�=�q��Ó�.:�*%#-�$�
����g��[L$u�M�Jf;Sނ��T�8x�wR�0l6�cBp���Ƀ&w�����F���rl'k�Y�}q Ic��E_ �Q��<�=Ȝ*�� R<֟��Ɏ!,�f��/���~M�}�³�tP����4�wk���%MC���nf�E,�|�B�,��p5s�#�t��_\�׾�I��Z�_�+og}��
��얓�%�2���e#|�!����H�:#�ˆJhZj���ob�oz!�{��7�;5�M�%%`���FA~7���kO�"cE5Z3��ǲ�1�B�V]����G�e�S]�G[�����{������o�H8$Qu�,�1���e��x��^�q?g,��C���������,�$�"y�a�H�I��,]s�X��Z>a8�B�����0*3�u��#BN��7����_x�x�c�ݜ��6jz����)s�˝�ȄMp����M�����������b0����`x����k#�6��y�C�"c�5�s��6�$�����̀#.<���X��� wX�~����QUcw��#�}j�g��g�D�	��:��&��������"R�ɕl[�
fOFRTiRշ9�-�k��w$�B���P"3\O��=92��� X�9%� {��*9����b���*�Cu�[M�L����"�x��2lP���#��DG&�H��0ұ�z��3X��s��ҩ�(���E�+KZ_��6kXlxVHYEB    4ea5    10c0j����Q���#Zl� �E�K��Gp1H��V�03��n^%̧�cZv�i��[{=f�m�n�����G�BR�1{C{T[��LM����]m/�XV���~����7{|��L*���_-@�ݽ7s+#%\vv6����F��Ǵ��ZYD�z��9"�>�o!m��~	�1=��kp�w^����<�9�2+뙓#}XJ�Q�"�
@إ��m�m�I/O�`@��kݍ��Ԅq�UE�N�^'6_�xV]3����K�g��4猹*⫂�w�����g�w����A�TJZ�f�Kh��8�l��C_9�F�����_���%�%触+����Jb�N+�[���D-���#o��j�Q2^�	�X�[W�9!Fٕ��?���~��2�6{�����t��qG��e��Ȓ�z�#8�Ќ�g���L.m�������_��!���mB��#��<o�UM��r��3y�����Ä���tIB�t��)�V=�=�1`4僎��f�P�D��3"�2wf�b�r	8H!��]�h�%�dV���J���
��&�0�k�;ST��X$�8�uu�	6��5�򪿰oX�
����n��F��/xU�;c����Et<Z�q<�;sEb�D7�lͥR��B�rMB��^��b2�|�t-S��xL:�+�d}�r����t<��VcgD�dU)���M(��\�\v�Ru\]iO$AS�R��6�/��`�7sw$���%{�I2���6CV�د�s��a����ˁ�rK%�P�jq���)�_d���$$>��a���bw��>�	S����I�"����4(�c>�'�=����8���f�]�1s$8 ��7�J�����l�r��Ӿa!�F3��G��(���G��B�mSi�VI��
N����֣:סz��"�@��ʜ��Y��u#��SY�$������!E�,����j��q�ɛ���m{&��)�(�U`�|c+����w}!�$���:|���8����Yٙ��V��E?�|�4�a���99G\����eD���e#���lMr���@�.�����DE3Ug�D���b���þP�s�\����-&��6��I�T�Ι���)q��R����Qp��T���G}�>�U5�pv:��)Bì)���B��J�;��x"�#~d׋4����w񧋴-sS>����i�h�/��}v�����(��Ӱ{+��X��qOE�'=)?!���W��S��،S�j���M�@"���©֑z�N�bKyz�;is9�2�@��ےгH6d��쮥�X \�*-4��1_��2S��A���\8��f��	~���4"��+@����$���밂�5P"����XmQ<ނ¦��O�`Z��KD��ֈ��R��50]�nf��0�x+d����=Ծ�:�<�'
��W�|d�m��Dv�@ϒ7g���K�t��w^��$L/�r7�G�}�'J~����&{�p�ʴ2�O��?ŻD}\C�P�ʖ�Y��ܶ�%q��^gIJ1�헏�mϤ�3��Y�V����GDp2%�W�=n_��gjo���g� ��fk�0�����s_�n�������В��k2}MwR�t��������d-��5��<������/�Ȧx����&�xg�G~��G̥y>�6��Ռ����s��� �	.��� _�U���K/�N����6-*�,�/ح�b�%o�,-����H�� y4�w]���b��8�U�fc� �8��7� }��ԁ'�C�sk
����\׋y�s�t5hP����ݍHa!W5��f�sХB��: ����R��O��Ëc�":�����f���1[��ϞT/j�]�iJ<���zH��#3���t�2}�%N6<���Ug{EL�+=Ut[s�0Uǰ�l"�ޯM�>.��S�wU�	�����Ӟ��V V�!ܑfhp3�rb2$p��16�P������-����Q�K(ذ���4|�;^��=y퉃��Ib'�ق��B1扝�-j�� ����
�/*��ᙞ�[�}S
���W}(�!�e�	�4�����������:me�|��y�v�d��܅���ğ�[.ȃ8�S���i��~��D�Ѧ�\15~��u����X��mC��ؿ���U��4�q<��Ë��}�X՛6�r�|�#�b$��ʐ����筞������$	�ű����Zx�1�__,՝�#��8eS���Ar�i�u������7J��iT10��I��i�g;ϲ �E�Bm2<B��g,T
@���[�x�=jjuI�1�_�B��p���Z�I�Ry���y�Sje�������
\ĉ��RU<���RM)�0$�!�<P�]�c�C��b�4p3�=1:�s:� k���E�1i�.���V��vb���v��(�"b��y���/ɘez��t�(5l�BȄ=�`�$R;�D��W�{�<|ˍ�ҡ�������T_�Hm��.�1�S_��p�'j���i�H��;E��e�����7�<��`'D�4��>!�5��.(p��s��c5���kͶ����(�d�	����9A�9��o�8����l�6��$O���IϠ�B*��HO�!���\��T�'��2�]p�^O����q��1%�Xkr�Ջr-�ڡ��3��%B
+��r��w!�VE�lT�g���8�����=���%���X�+s���K�o�G&(�����.2���B`6݂�����+i>R����ݣ	�΁����:��b� ��=�ID&�3���h�W-ZMkP����!�$�]�x��+�<��'Q� �m�$v�ƚ?Z�¬󍤦�ŋ���~m2�����5�[/703���ĥ��R���7��~�-���ѧw/���#�e�X� ���"ؗ<�>(w��(�����y��j�u���D��V�cɕ�K�n9c�v�Z�_�w�K�>Kz�7��o.���#��(Z�U��^�'7�U������ .���Z>��;�o'�Üpu�7x(k��?��7<o��^a��=P�Q�߀��j���t��d��E����y;󐠑�!r|�'6��RҮ�7]q�
f/�Ke��΋(*�"��Nc�=�&��A0QZ�h�R�E�iJKf���.�ר+���!�>��U�}PG	�إ*	��� ",�lԷ@i��j��	(��I��*�7[;<��D�k_D�^�Vs�ڽ|w(�8�kߡ��1Ջk9�Y�Į��Y!v��\���a��5,0 P�4��jȱ�f��f���Iʭ.Փ��L�Y`˾�=�ߋѷ2Qb$��i�����/�?j�����f�$[��3�x�T�ɓ�h��iV���[��vx�4tg�p�@�5���
r�:���7ֲv� ��\eb��x���/�M�<�nI�A2y�,�-� �Q�]����~=�D����+f�sp�r;5�=���c?�c�;��m�g�>r�hvUAir�����7�D<�]���:�:�S��j���U�F�B�d �� [2��_Q���$�)�Z=Q���HLU *��Z;�*�RK�qI�M��N�V���ȶS(�p�H頁�ׂ�*JD�}`u�2�l�̇v��K{G�Sϒ��e��>����<�z�xn�����C�C�g�2va7a�mֹ����Oq{(����(��&Ha7�d����ӎ�<�5�?aoo!�W̧o��ĂRQ��+3�br�5k�a�>C�� Iy ��{�KԤ���~����68����4m��7U�_n-%
H����?թL^&����ht�M�M�����څ��/yh�����a>
e����&�Ԩt|�����L자2ĉ��N.g<��3u�I'� 9o�JPB��kE����v)ar8�nm� �و:�K��ӗ�`�wa-0�V1U;Ǖۉ�ϛj�D��uq:�T�>w'6U��E2g�r#�?� �O���m����f�Ȼ-~�[�i4�ͱ$��uw0q~�� �#5�Qh��T��[ih���������Sj ����3�n}�k�����=-�8��&$h$�k\��]ƺ�kPpi��^_�%͞�i��`��jcc��������濄��9Bg��x��g��Iu�@�����@�2p=Ig@x�G�fz���������Ӏ����T/A׏l��ٚ��.��E���gUaA��&�mi�;���GrH�l'�+