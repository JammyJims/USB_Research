XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���&DF���S�5�R�����)�ӿ�gR6�e���J��q[7_����m�0%X�,a �0�뎫��k�~ڶ�@�J��m��!��d�)6BQ��E*ɵ�f�JX��Ŵ�Nl��{�C�]��}U�Y�L(kן	5����IXeG��t�C��> ���uN������Li]"��)��� �9XH #Un+7�ׯ�oF��և���!@�Z'��J�.��4~�yՏ}>���KcA��$�M���w�<�k�t*��A���>F�R;i��}�;��F�n���w�����ep���w�n�уï���
y�aV;�Q|��z���D��W��@K�?��e�a:�*�����[ @3ͣtC�vY�t�T'J�&%F�dw��*�4o��?X/[;���8���Z��ta���U9&&8N J ���> ��q�ԌdF���t���qGzL�{h�L�&^%��ș��F���b$�(�,��� �C_d����U��� �������>T��vF���k���F����G�%*呸���=��H:�9��d���i��������5Ba�D?_�B�&�/��d?u��
�i$#M�A3A�N�~O���M,�0qj��	'� �h�O���U�n{�*�Y�1ٞ\SJ���׍�R�8��=\�y�ĥX"�����T`��H���f��4x�������nV�;9wR�8J'��^/�οK�"��ep�9�q�������/R�G]0͔436�V�DXlxVHYEB    5765    1330g�����8���<�I	_J�Y-˗��a�3��-*��X�L��d��(�,��V��<G�I���&w����h��do������}hK$#���.�-�{�j�#a���٥0�Ont�Cf��`��=u+��YZ��%�j��E�� ����M�`�+�X%���g��l��5�p&B����7�n_��C���:ʑ�?p}��CM�A�e�9����K0A��[z3��Zm$%�5Ik�ze�B�fWk%��({�@������&YA�G��s.�o�/3�SE�b\Z�|��}����G�O�x�u�7�%Զ~[U�f|����v���q�e�.�bj���s���]O����@�NY6@��z	�n �O�ts!�B:���;?g}ZCq�w��1���e�����s�b��b)8��'��?�\Vw�)N��s8��s�Ķ�#r׫O�-����n�:�y=ęϘī+��KHh��@
(:��->�NF+H��>"���iGa7�,���ݡ@��.�w��7���9��s!8Fĳe?HD��^_\fXQc��*�V�:rF��������D!��r�n2 �a�(<�DO����kB0�7�{E�%_V ��d��=�y�R�k��H�4��F��[� ���)�������L%~e1��� &�/6|~n��K]9���dZWk���n[��l_���Fi�ȓbTPoB�K�Qv/>���
K��q]���/Xw&��(����j�;6q�<8�G��9�SH�>�8��,
1�Q��X�c��P-y�2�ս}�u�3�ڗ��bd<��/��p�'m4:�53�k�롺����=��9b��"�f�A�Zgu=$EG{���{�D��;�����Sh��[���X�5?��}֔"%%+!�<��O	^Mq�0�	��(����������	�o4t��q���֢�V���Pڮ�@]/v��IA
�`0��A��K�T�%�(2t��@�!R��G����=5��juP�*^��>�1nix1�TaV�(��~1Tf��wm�gT�6]"�Wǚ��Yf]F)_�˱���t�{�"q�?��s���F�RP�\��q����S�5{��q�*&�<z��[0�q��D���ױށg�^�
q�>v�� %��"��l��D�?yi*����O�>#r�/����
����,��n�1��ǃ��W��?�[�e�y+��w�L����1&w *z�L Ǳ�3$^AF�������p�l{�*/��2N�p��~X�g��@�	�T�F��a��_}݊pG�����:�M#f����������[�l�M� u�"�n� 0�n����zT�ӯ
�U`c�Vc��8*8��^�mi7%��TK�`��{�x�@}��!v�O��@=�C�KuU�:��{p�����4/�x���'����Q\�}�b���>�2{�Gͳ�@� BH�/��q��2:8.���������L�Ҁj�c�]�)H�ybc(�߼Ai��c�)���E�|+q�3�1�Ls+�p!.�@�D۩���d��T���`ו��K���ݺ��k���Ƽ�c�����<�sM��#$O�[����5�J�Z���~����1�F��1=�7Ǌ�_Աw�|9��[g��=��p��wޖ���,n����n���?�}.Q�R�IX3�%��y�eh�V�F)���؞ؔ�ѶWd(3yg��N��%>�~R#��I.�(�;Q'-
�gYU� #��J���c'�[���:ǉφ��0R9������r]	yk4� <«#��H tAP�n@�MB�.�0��I(X���41=�'B�rNНXu�S���}��z��2ÚJ���Ě��Y�I�/E ~.j��1��0��,��)�"=�ޗ�D�i~�GI�-e��=s?b�TyL�
���^�a�5k��RD�����-^��A];Ff}�2^(��]{�jK�7x'�ST��vj���d,��}���_�˓��EW�&m�%�}���D�v��!H���q~]�˃g��Z��/�2`�pm�QKi�%��+�T�ej���M��p�gQG �!�шP�ϟqc��V����yqM���>s��m��fNu��K*�Jc��)\�cTlT����cN�t��]���78(t�d2}ë9�	%1�^��~��SM��+��K��o�o��nߺ�{�z�s��o�0���^��d ��)�Wg'�{��h��gs���p5_��لGE	�$���4�����p�C��>���N �,�LW�{^ó�������7s"C �Y�ݩ��/SR-�-_�Z�5<�5��J�8�GI�f񗃻���S����n��w�o�����%bd�}��@9��Ͻ��9�V�fPm�����*xa��HUe��h%)h��(7�g�$���el���o�U-�?�v�n��1��#�4�aM�A�=g�$e�gl���HA�yr�輩	,��5ϔnIN�eR��������Q�p�T7؁�І�G:�;���^��pT���(����~k��zZ0�M,����w�>��V�e��%��HJ����'w^�)�8F�T":ٶ���KǙ'����p>Ny��]@���H�SՉ�7����\�i*�A�6���~��Ŋ��G��%E�t�t���
�OI�;4P�SW������&+�j$����*B �|j^�M���aJ8���%{*h 0�Yj�o�	5dDx� �j(߀G�]�p�0Z�6Qs�5�A���Pn�l]�3���)������s�-XI/�ڹ����"�������
,9��_��3aC@�F��j��O����>ÄB΂b�����e�Z���GG]Ӂw���N��1G	�=i7R��6s_Q�Dw�&��������Nݏ��~���υ���]'G�kh|o��cе?~�%��W�P��F֤�r�ĒY�P��*Dp	�JԼ�ʚE��,F��%�&.u�u�̶����Rj��4r��d�=fh�Uw��e�Ҫ99ؕ|63]U�����&7����{J��Y�3�s?���X���əϋ�w�V@��@�=�G�p,� =�c��D�a��5r�����B4H��-������
�8;w�?���HZ2�?9h�Yg��g`Հ)y��"Lu���Ct����$��R�\X��ct���nd(���\~�7Υ��; r%;����P��-1)�^s�g�ǓX�m���a�9�̶Nq�mS'�-�m�Dg~];L3�����j����I�J�bݨ��G���[퍓CtE�6�_!�6�>^�J\�0��ͪ.*�!f�*�Ԕ쾤��0 M��!]V����i`�����6yT9p��a�t�z����H�Mx.���
)T�Ҿ���M�(}*q�qOܖ����t��f>��	�M�,�k������sdux8��s�)D˽I�}� e�c\u�3�e,�A@�T��U▆� u"�|�&<����/Y����c7
\��M�,��yτxM�c8�	�=�>�b��p�y)���~"���'�J��jx')��ѿTl�e��g8(?�ˑ�{(�ꩢ�|�p'A���`��Bf��[]mL����T�ue��
�$c0�N£���^��ų�ќD��(��W�A��ľ�1aBW�uk#�3�:"�$���(��Q�4�YrK��B�|S"�^Ka��|������z�@Q���l�x���½����>�%�ǘ����5W�AH�m�!Q�4%�ENr.����E�������m'o�gY�r&Kn�|�i:Tr�|w��;R�c��|��������Γ[���*%]�a|�L��H�vy�2�����PgR����bU\�5|����ݟ�"�
�c�Zg���G@��	@�_ֶqx�y����,�c���ː��&b.�P��:�K鍓��^��s�3}8(�V��#���ú[`�A���L�k��R��SeJ1d]p�O&l�eף���l�PP���!~]�;��Mq��U���1�4�X����,4�1�<5��';�4"��U->2�^aז�M)MӾ���.�	��k߲Ěo�}�/�3�=�r7���8BU��-�}������7:ᥢ�9h�3p�'��׉C�"�A���
.�;��e�}P� J���c���*��l�Tڦ/;���~�P�T"�`�8�<PdyX�~����ցV������)S�2끺�Ϛ�N"�\��{��"���JG��K�^nO��A�/��]ulP���2���k���A9� ��*=�J�#�6!⓿y��z0m2Ӡ�oB�̬�9+�;v�ҳ����5�m֞�Y̤+��`��N�����Ăe��Fw�4ɐ��6t����i�t�y-����c�1��[�ǅ
X����dA܂݅�����}�p�l�/%<_���I��3�U�(]@��Tv�td��:!bW��-v$�e�.�@�	w�m��ǽI��}�#7��<u���)��{]i��$O�����"~:h��GW&���Y�d:�FVf�iu�&�_moݲ����y�})���A�xAE��=�I�����:�4E��tb�g07�4�a��U�[�_�a2��F���z��O��u�U{N��E�3󿜲����n�n�]�ی ��C6�ѻ�]l�7�-�t����<S�� �U�@!�Т�t��9�DSU~�s��p:8:���P��X�	��Y+#ѓ�Qޗ�p�zTv+))#&(��ǩ��4���֥�Z�٩��{���s�	>����Bb�T��'�V,+�gu}������u0�0<��)��?�O���,9`!ׂ͊k�	�M>h�S6�����¶�WA���|4�p�9)zN{E�r��