XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����_���˰�(��b��x����a�WD���q.:�(����~�O4b�͗9O���$�g%�������Up�0�� �"a+�� P�f0m�Cބ���z�[[�Rӟ�"�ŧV���H���%J#)�6��@ �9�a�V����{�.� ����Z����E��,�1��t.-�8W�m0��-����+T�]X�"Ü71˸?a��hL�c��Z^���BR����>,���k��A�̠�I��i�x"�ɡ�����Z��C�B�#+�$������J�8Ty	���.���b|�rP������Y��"���
[��o�d�eh5�"t�B�U\���}��\�ra*-5�>�5"��Ԭv�΀71D:����ՓX�&�C1�<~X�
��uߔn����<�V��A���J�OzP���w� ���1H�-^��+	7dU1o�VR���f��IB�p� �,���A�b�;U���H���`�X���F"���3�Q#��	An'��ϵ�b�A����ƑAf��Ǳ�+Ni�P�	��|�4-���!���^_���R[��]���H�q�Қ���ֺ�ϕ����0=r�<�6Y��5�!H#Th0�)��WH���oL��,&�����NPU������+��/WGL1[]�����KY2�k7|��\��(�wz+�Ze`uÉ�I�K�_�i�|��H���t�
��B �`�	�^v����7��VG�O����cڍ���uʕ�z�o��XlxVHYEB    ab4d    1f30��������л�˧&�?0qK?Q���/8ڑ�0|j��"�'�\Ҥ^�����AH{ 
�'����������-�ޞН����(��E+�4'c������AS���y}R�F˝A���Y�e�r��dcI~j�&R
?M���t��s~Q�m�&��[`�;����nv*��O:�\��%�Cؤ�kdM���{Dt�I�u5�M��e1D�i.l��H�V8�6�,�q8�f+M���Rl�]�}���a5oR�l� �f����k%�\���lE��)�[3	�;֯ �P�!Ӕ�F�8bم�j�m2��Gf�/7JZm�B2Mx}5�`���k���KK�8n��7�.�[��d<��":3�'fdQr��|y����PPJݺ�Z2��.�k���&��̃%�ʗ�`wD�mf�<A_6"F�fʙ�doArE�C�=��h�̦�7�i�9>G�����aB[u����"�?ҡ��'�d��Ǭˬ��1C��*^흂L������<��<�ڑѸ�a$���6߮ՇH�szO����܉�0�<�z'fy�����ZM��nN��^��rl&Ƚ/b���l&y�7�����2�\����欻�����X�L�.24�q*C@�m�I�k�q��T����'%�.1�[�%����0�S���XD0�������-#��t&
�̅���:� LzYR)hR���K�b<�]ْpO�Dv ��|VSh*F(�����
#+"��çc���g2AP(�L�X�	e�ֆ^x�Mb�2�q�2�w=�B��0��9F�@l+2k�R��ȷ�c�B5=�.���pkq�6�*=�̿�eaM=-�g�i� $��i��-�rR����Y��,��LBy)߀�X+���9.�5l�5$m=?���P���j���o�qѪ�Ɗ�4*�?����&R�5e~����Y����.��8z(��r��o{L���O�3xAɝٶ�@>S3i��ק���sv�OXqv�$�()tR��%���+�T���*�P	iCK���P�()z�J��Զ���A,أ#���܁����Ɠ)j�TE_-�'��Cs��U]�[�oF�S��}j
�5��
Ǣ�V+�pTdG�IX#�80�D��t�(��{`qц^#���fQ�~��%HP�L`iڡ��@����"p0C���g�Y�bSe�ȫ��tqAޱx�*Zh�N��L6����
Тmy���]WB_��&h5
�q�:A�@��14qa爭��(Ϊl`��+�&&.��ǚK�%XB*�BJ1��i�%����:?r����6=�}�f���!p��߳�6�T��_�FQ}̪�����Ft�|13�ef6�u*�!Y?&B�	ڟ���c���Z�חî�����,�QD߈j��[��f;q/,_"n*g���I^�ʱ\%����x�?U_9�#����3�,���=ta�_�� SɷK���!����f}x8��!y�$a6��מ�c�3]+��Fy!���Lr���33-��������o�9
��FBߎ�j�b�I��3���x��	��~��EK�sn�?���l��p��ʶ���Wm%�ee �*.�u�7�K{��5j�3ca{�V�u��F��Jd���iX٫���<�g�_m�7٤/����s@Q�Rks��RE.�H820�����B����Y.��l�t�0�$�J�����"<~;�q0��MRޮ���tY	�e�\'��Y�l��\���vu������2�ðF����V6�2��°��1��d�ni;��wFw�s�f�>�=���a�pdѡ��.W�d�=#}/����"���DS �������Ev�Wgl��H��랟����ZpC��xOȢ��g��,\ʦw��Y�A��Y��0%H �I����_�M�׭�(��&zi�~̴L�ϱ����suڸA�{����$I��D#7�����.m6v�K�*'`.	a���6�fȂFx �՜���Jf�c-��#� �3���Q#j��F]��Ey7���?�k��aJ;�ڣ[��Q)�V�㌑���,�?O���f�:;�,�5���OgT���t���c����8��KC�P���lHP�9�m*�y��nVބ�J��4�H�_��1�f ����Ѽ�W������b��t��~��1:-�>��l��VS>}��[}S�>�?u?F��FV�>ض4E������Ļ�'��3����<?��rp#%����u
�禋�7ѷ�)�/I?|���ɨ:5W�Ӓ��	,�	7��o!ȸ{e�6�r�kÎht�+�o���Wz� �)	`�:F�kj=Ԗ�FwDӇّڙ�da�BZ�)S:�a���ȫ}�_-�:)5������e�l��3ҳ젺L٫��>�ܶ�]�SS7;�|,�����(YW��oBz5��
-�6�.�� I��:�g�	R�"��X�[��C�ޝ�-FO��,�>�1��+seq��]w�0L��J���r��B�=�AI>�]�0u��BG���g:J��#���V+D��H�9vMB�5���"�,����z�O���m{�\*�����t�&�Έ��Vʙ	��w@O�%G{MT��]��I5�M��&o��f��dػ�gCN"�E�� �B ��%3�j�.�5�K��t��zwv��<��8O;���C�O��d��;��)~u��\�n��
�8�M��t��B�*��SB�y����52
����
&���b5��}m!{���V%�WE�S�	~�E[��\����l�+ gMf�h��U�,������L�"5N��XB����&�Iduf����U�jlf�y����c����_�7��L��E�#���Vd	�(��k�)<a��V���1�dc��a��3!�Ih	��'ۚ��%H�e�(O���53$4����J�P ^���uY��!�c�8������QH��"}����wc�[9Q٪�5�d�"��"�o���jFP��� �A����q��@]�J"��_�-�^��6~�y�� +�60$\m���UN���l��ٶDp�u�ɒAM�����EW	�~m)g.�6,(ŞV�b���O�(��.V�/�X�8Ja��j=�f�HC�I1J�^~=��U��W�{�tB�uw햀i}��2ѡjj�t�}�"�ǞJ����y'��wC(�}nV���H`�j~x�6P��7Ut"�R�7�����0H�a��N�[�����zW9��%�=S�g��w�$�d2���I�� �-[!as��. iL"�k�Sφ�	�@����AYBO�?����k�ۢ��{iD�apxy�z�b��~�1a~����QXf�aHP
Dx����dO�$�Z��)?q�]7'��<����/oR�{_/���+t��Q���й�� ���_�T��DLfFE��$�D���TWY�����>����0����t�v�(��R�"r!pɆ_&$�}24	$u�_w1ޫ uY��!50���8��i�cDO�F��Ύb�� <�ȿ���z�,�#��P����J���sw>�����+_Hۀנ�Il������mr�}G?)�*:����_�ٍ?��3z ��6���Y��9�IB�dO�e߿x���E"L�J���0�:?�k#5<Q(審児_V�x���CJ�ޚd7~W����;u�U�k��$��FoZp�5k�IRQ&k�3��k��s�o����^�8��i2�a,� ?}n�l��y�x����_N�(�j:Xb
�y�E-��B[���.z��hW?���Eyp��ib���,�?��'����ɇm�o;���*K�,Iչԅ۝IH���Mh�#��k�$�B��HSv'�\R"]�%����.�få��J�>���GMv�x#� �����ì\��A!�Md���\�86���Yi^��q+�h0�+K</k��*��2?TZ�r��б�<&�#�5Zp�M=�ڿ�9LE��x%�\�m�T�c���^����������]�fbh�	!���	�'�P�S�E��j|��^��{�D!��I�=��(�#����n������v��9-�	��*kM-�E:�N+�a}��ۯ��o����Y.�3.f�Ҏ�3cX]�,	C��E���3Rd����������4:�腗M���E���\	`*��e�����n[�J&c6�����u��^�n!0{�.��a�?���W��G�bv]

R�W$[嬻6L���k��\z��jga������0�x�`�APo��k���O6_u�9��zJu�_~O��P����۞o�Kt�k�U\�������"Zn��!�V�կ`m����i��*�$T�6����߶���J�D�wG���,��$�D�r��ï� �;*_�p���ڲ/��3�|ǅq�5�c.+T'd��,�Z��Kn�<F��j[�z�`�E���w��DU�{n���N�|���ߜ��{	.�]�*v���.n�w?^�!������"��@��	�FY�]ٯ�e���U*/�����q���'�?LW�������h82!jD`�O��n��1Qh��r~�??gA�`��y��s�lg�~u�!q;��3UjC|��k�"��b�xum9.�cAۤĥ�jy��%�)'�V/�p�)�<����;1����T�jk�+��~�-Y������Z���؂@+�JQ6�x�t0�܃����"`�C u�Xʡ_�ZcFj�v�r�T�������2J
�Y'F���\z�C
�f���Ѐ���ញ�Q5W��T��$E:�2 $և��Ppb�{�7���-/��xe�BO}�y�BbLl�/�-��}�[����ԙ�ew���;5;�����~�g���ii��֛:��m�䡧";i~���ȡ�Jl��w����Èd�[�EMB:Gl�*m	�����aZ��6_F���J�Ռ`�*T�5�2�q�E11�	X�B���?$�*	�ى)���s�5V�6s�3���6�X�ds���<e�v������^���.q����녷�'@*���$Y���Q.���A��ܼ�b�0��M4prX=���dLWZPi;ΣtGd��v	���s��$��LT��D[�ʄ5�H��N�-�ļ�򉰭�:=�<y7���|Z���[��yF7��z��}�l�� Qjs���*�;�����io�р�D�&�&���9 ���ً��^¦��j[���w��〿]��N�ט`h����OY~j'� ��J2����t���ʗ���ymR����EX0y�8�	��zU]�$�U�;�"��/�-�9��Sʢo�P��$/����Ϙ/9Z�u���3qv����'�c���q�w�9�n�A��^��F�ժ�Z>�2K8�(�n���	�0�&�:��c*<քsI>����3��D�r�'w��X�1��yz`B�sS&a8.����){��&�hgß0�]e<�)*���q�,Dm�9K\"��!�w]������Pמ�J�no�u+_mc"�2�+�0s$)sD��a�ϩm?�H�`D�Y'w7�l���W>�I���5%;�"���M�� x�<;��"���^�O7��4ee���䧋�]�ԙkZ�qآ�7�A�//F���a|��v���^�?�o��0'-4��jI|�0��nq�s$����q�?�Nn��K%�2ɪ�^��ϐ�d������AQ.�QkalH)�����0�d�~j�q`����I-dn��R��E!���p�/Ā�/�l�p׋�꼊�yI�*��5������tUvd�]�T���sY�,�/$
=�����(�06�0),������O��<<2���u��ZH�v����sz#[X�<���i�/�4Oݨ{˅�"��1v��Ċ����옟U�%���N��=ч0􉇏c���)�ɒd��:j��y��X�u����3[���������B5��j�b������pt��������~�+o���F���Z��&��Z��	��/� .��n�b���@L��^P�4�S'�88�}N;��ݎ$A�?0_����J����J���%ҿp�/��-�W�?Z�	��,Jr�n,9���w1\�&/���nD��`b�M1Ѫ���qh�5W	0!�� 1*��3a�g���=��Et�2ӂ�՚���ͅf�������s!@�#%��,ҕ�t8�C)so]1�8�'b�kQ~�����	�2�Q����U�Y�Ⲧ4����Ĺ��,���+�)YW�5�^���4��B7�X˼/H-�΍9��j/��������X;jd̴,@[v:D7|ekq�"۽�$j
������3N��B� �C���AD\�� ��.e�4�4�մao>F�v(���i���]x\�*����`THmr�E?v]/1}!�5�C���	��3B��=���x,V2��s�*Jo2�ݱ`B!z�Ji�y�&D�mi�L���ʱ�K��H�mz5����4��G�>�)�v|=,�6����v�]��l��R���s�v�b�CE3;0��(>=����2�h�~u�3���G欇3X�@�Ž���x�e���T�/�;�)Q�u��M5 ���A0�������d�z6��;��$��>q�n�Yt���Q��[��#l�w�"�r��K�tl�Ci�|\[5��t0d�w���$jܓ��e����渝���L
iGp�Gp:�_�A�WW�\!=R�y����w���C#�x(OpwT�\FpI`�@�� 'ɱ���n0�*�����r5��}]y�ɻkFU��l��m�M̑�H�r�^O�Q�"Sq@%�'�W���e�k�� p�v�C!]��Z��-�%�g�����!Pd=��ˉ!�����[w!���mNP�K� �0�\g��U`JПC��G�D�ym#�c�O9֊L#�%�.6O�s�����[�}�0`��$�izm�ܐv��K�C�Ă$��Z�qZR�}ۮ�r}��\g�i{ۜ�?;Kץ�ۊ���o;hHs��уn��|&u����4K��>��՞�9Or�C�.w���6B�N���0�=�Nc$�6���G�I�o�m�s���u�z^-�9o��	�צڻ���%�`��С")�{��Ĳ�,	�O��� [Fj�v�b0e��`�e�/*�y�s�B�;�\1��'B�ߟ����RVC�j@�/f3�Z�L��l/!�?(������	�R��2���ŷ��QJ{63B&Ԩ�/�>�w���YA5~*�n�hBʕܑ��QW�g]F'W3>4iгom�Q�O^�Z�TJM]1E��i;p]� �T�C��9R���V�s���o`)�aQ�d�9܃�r@���#z��Ł�� u�tg��O�O\����lyj~&ϓ��]X9�U�rBn�H=���W:�ȇ�*.ST���p�Ք��\��=���An������h����ޤ��П��0xZ�9��J~��(Ӿ\<���`��
����\/�U���H����:�ƈH���dr�/|��5J���߻N5�msw4|�dT��8� ������GJ�Y���̊���4��:Zxmn��W�S�����g�]'��MEi"u�������#]J^�77[��P�|K|�}\7F��IK�HǨ��Wi��~h�uO8J�q<��eo5�����՜�ҞI������Q�X}��4�����['V��z���t������v{���VF�h�'f������_K�_�q�~c��dU��<�DD��lk�_�@���(�G���Š#i���n��`(�\���9��6q(�4�Q�$6�ɩ(ޤ�*�@�n�6��t�zTuz�$RE\���O�J #�J, �e0��cx�lje`vA|�@���c�g��L�2)D�!�B"NM}^/��ª�ԙ��2�e��f���ݏ�