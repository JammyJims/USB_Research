XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#P�]{������e�þ�̚ƺ��I"�ĺ���7n\��?sj���פ#��X�]�����÷f-@-��k��J����x�h�GA)&�5id�U��x����y�[MS��|,�N��%�K�����>�|�g?;~���x����W��Jq�	���IF��)ٰ�e.r���(<��;�7b�L�+~U�F?tc`��3�fS�pf���0e��`�$c�m�*�7�r B�8tq8K�6s�r{��{>�r���$!2#+��dL���VT2��M��{��N�7dv��&�����|�5Ūhn�2�K_Aj8%��v���\RJ�oD?�%�4��`����[l��LM�q[��:~�t��\��6Ԕ�f,�zS>�w�рb�Dw��pFH{�K�Q�Jg�!��H!�p.
t�ӊ���&oη'��`�]	�qsX1q�a�n'���z%��4[*���3o2}<Hd��h~� I���L��	v�K�Ҍ��E��k�/��9�H��?�G���v�5ȃ�
�pP�G�;��}�[�㢚	����=
 �ѭ9�6��n����-��ͅv�%�!�	����� �`%���20�h�ޱ�eG�|m>�l�E�u@з�Gagia��#�,2M�W��^�Xk���<#���\�f�J������Y�[�N��]��{�;5�[�It^=Cd�L:ۋ~�س�����Q����|kx����fG�W��5*���W�L��ܭ�_NF!�9�9j��k`�TH}m�5�XlxVHYEB    1ab5     7d0F���L�8=�$W�X����/�Ф�v���7}M;o��A���k#v�N�G�������Q��\�*�P�W�p�Lm�,(��\`��'�ڢ��4��g8���̽�%^��.���r�0�{�ӆ+l��($ə�5'�)��d��~����!Rp%mwهE#�E�|J���c� v6QCV�bQ��Nhu���Wl�;d:�z��v���U[j_6l�#�M�?��ZG�I�z�t���C����tn���m�c�`�}_-wc���X.^�ߜ�O���ym�U��@��h/5	�C{�-�n���WM�qbz���h��[�w3d^���a*n=̧&��5	�����Y�%D��7l�r�
�؋@bj@o�����U��R�#�5
ϕ�yT§�T�� \L��_�foX�p���C#>��
���ê���/��U�UE�a̾�ɫ0U�z_���x,��tSe��{Fl��+mإ�	�A��9ۖQ�N��W|��S(�Xi��w`Ǔίb�������EV�^���[�J�������d{��<Rs{�i-LZy�캘���9�@/h�xQpD��1��mT;=�(j����~L8є���h;�%��k:�)�&�)�g�&���X� u��g��sb>��̯�cF�!1���. ?z��L��TĚ@mG+��<+��|*���G�Je�uBY��:O"C��E]�Ne���ԑ�JNצ���oW���wnd#��{��$-��@���eN��ǜ��8�r��}6)X�90~����l��_��F��:���Ժ�rMȎ����=^�&0K�.���,p��,q���4s�u�a�3ͷ�<%������17ܫ6��cs�Q�J5��"L{���0P}&�n�Tp�>�z�Ĩ�4V�ߒ��zŶ�1tS*���y�!��^�&�aQ�C㥅�b�=i��*
̙���S!w�%ق���x�pX�
i�?Ʌ�2̨$iR��;���X� ;����<����sP�b)\�1ƌ[�=`�Q������|�k�"�;��z+A̢d�oh2������ﴋ�:�| �L7Ч������j>�;�������^}��ˍF!���Q}��4�K��KX��y =!���j���As�W�=w|c�� :w:,��Y��eЊ*�u�%Q_��.��(V�HT@�"W�ԇ�H�'�jnL��:��G�@ġpj�d�����f�1(�%&z?�xO��\:�씘>��J.���Q�r�e�j����:�E*P��o�hD���=��S�n��ա?]��Z�$�J�7a��qH\�i�}9�A>�Y̻�9jΚ�7x�[�X
�M�D�U-ud�9<��@��K���jw����R��M�`}'��|Z^(n����h�t��O� ��p?L�Ӭ�`���Z�qrP���h�]ü W=�C�.�.\�$�6�3�Ly����&eJ���"'.k���Dm-�ߴ�O.dY}���u�������LxTS���5�o�o*9�.�����t���9ӻ��т�)l��a�=� s,��H]�p��'���=��o���f�Z�Z�Y�!-�+*�רd���d�BE�4�C�����#��<~�DB��n;g؆����,WԎ�{$
��!?�7���1.���r�R�EK͕y����ȷ���ݲ8��x�U�J��1]On>��?����R7Չ�>�<��{_4z��`+u����stח�kd���I�^! �*��z/ہ ������oM�!<��pj��r��9����=�y����J�ߪ�%��`!���֗�������mhY*%���͐�@W��/�|�^"����ڃi�����ϳ54��%��g�U�%#=P_xm{뚕�����9偡�Vm
��?�p�U.�)�t���DG<'7�gʪ�CM�<��b=1�rۋ��ƶH?����"l��3������X*8�|d�\ƴp�6�