XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Xon���Tr�?hs~{��$!��_�o�(h��K(�_��sf1"�ƭ��}6$͓tӟۉ�Q����O�����4:�T���e�zC0W���x�c(�˺�3R���~1��a��"#��*I:�!���g�M�"�M���2�mp�����g� n�vE���ǃƃ���n���4q{�t��HYB4=����zMn[�7��#����`�~4���!	 5��l���a�8�N�B��s�6����ȏ~��ֻ���oܕxǉ� 4�e��_�|��i�O�ID�`�e\�(	��V�w����&ϲ({��!I�t��h��z��.�E�<e��"��p��.h�M�� )?��(>���az���$����S�J�|���2;kd)ÜP��K�d���a71��r�N���Y�!z��H�[jLiD��B�1y��i����"�;]�<�d�z�C3�a�%l�����p!�ˇ����0�B#��˟��.���JNH�:����>@&��1CJJ�SF�1�L$��[ޥ\ur����7��@�L��ʄ �����4ኬ�0^g�v�����8�e��U:%���_08%i�0ݠ�q�!�Z�h����l&���f�|�$^{4�F�O��Vp�R���EH�oi7�~���G���������G����ά{�V�B���^�.�_���������
1��� �s�J�z�E��A�禹���w�e�8�������;��v�Kf^��-��XlxVHYEB    1ff3     b20Q�j�ܧKv���Ma��ګ����`�31Q����t=�?;���q!��Z�p���+���7���6w�Jr*m	s�C���!P�o,֢�t�����nD� )|��F�{X!���~�qY�:]����\���p^��6�}���IX:�%��g2����A|��ԇχ[��	�����RS�CP�`�Vw��H��C�Ѵ��T��A���J��.�Ɉ|{����45��4�Q7�P����I����I_W�ϼ0k.�?��Sj��ѿ�
-e�w�l��BI3�g0<3x��
�8�{�H��C��� i���`;�G�$F��4a����N\��kP���� 7�<�`�_��Wf�˸�ݾ.
�����I���䭯���q:mTs�ڤ�r������'ͪ@/��[	S����[E�L]��^��e�e4���H�E�*R��>?�Ϲ�]��YV|���9��#pY�����g��©c
��ߋr�.h	�Kf�+9!;@rQ5�+����W���X������%s�ZEv��)B���LJ"VM���ãn�'S# �����v��ĺӪ�5*�k	��'�6�-V���(?�8k59lFJ����%�>��	�%\�/��y�io�Y���c(��'��5���ͷV��K�(�i�Miϛb�*����M\aH�D{��"�Ȝ�������A�:�*7��.��e�a�u��]b
��p��|;lW�_o���(�k`�����\yd�X4?
���� oZ�����?�c��n���:~�a�l��g���z��`FЙ,8�� h�at
gx�;+fp�k��s圼�\��4IŴڦ٨:�%&�0�7V��pX��e^4e:���1��K>�����)[i��5l}�z"[!3���U���d�~��9���=A�B��>&E�W���T��M�!0Y��(i�@�(��u�(_j�÷��g&��`zO�!Z�S���/~��"�QH]�9��#�����u�R�p���\d����&����B%��.��L���Coې88`�t{	@��i�� /[��E�v�;��=��ϑ4��X�>X�i��ݍ��?"��ҐV�sd�d	|5)g���d/�M�#��5�
����n�!"&��;J���r��,Gc�Ph'��7CL���ep&�!�+hD��[�Jyb"	9�Gwk�ұP��(��B�p�P�!X��<���ĕͶ�fuo1g��D�4��`3�E6�۱J��53ԐU��������b�5�nx� �7���8�?=���R#/lMf�w����wƜ��¬��B�]��WkH�����%���Q{;�N�~'����S��E���cv8౜{{
�s��@�qouS��Bk�g�"߂=E�N��CW՟b{m%8�Mk=1���5]�D'0c�9V���{3�AI�'y���p��M-M�H�.�H����\���C�F�2O4�98]���+HR��φ�p|��\lŴ3"u��:EqT��u�Y M��|6m��J�i��B�_�ќH��<�&.��B�W8%ty��s��u*����l����ĕp�Ѥ}����pGY��V�|k��G
�lv�؏6�^�%(o�hiN�2���)*nX�9!���.���m���a���ʬgZ��F|G��a@�б���}�uۂ"�4e���)��o��]���n$��,�G���s���.�P㪃s}�e��F����A!�cĢ��"�5*�ل�łYݩ(p�MG����Ԯ���A������	�����E�S�8@�,PG;����i����_딁d�9�q�G�&�D-���㩹�]���
�(���eɕ����[�`��,�4Q8.Y��͞Q�5(ᴀ����Z�ψ�?9ܠ�
���R�ܡ��IԺ}�j��|�v5�=��(�w�Z���3����M�C>�t���,�w|#o��Sԛ��| ]l�_`C���z��1Ch�q�w������`$�Y�gM��9���A���I/f�_�����]۩��wr�n��<�J��Y�˄��o?E������ �d�s{�8HUJt�t(�Р�VP ��B&5���ufkm�����eoI�����X�|�F͐ӟ�}�{�.��ϥ��_��%��%'��JO�,L�M�ր��"�n��i��{���nd���wY���(����d���D�G�	+�ё|̖�/��z��
>�k�B� `S��n�SJV#z��G��'�ȴkk�W|�M��clԉa3���T�E��(�X��%pUp'�m�#i[����g��W���qϮQ�ͧVnU�z���q�Qp�,=�bҨ?u�[�zy>Gv�r�9PN�&�q�%�Hi2(���T[�B�|�=������ltZ�À[��������=
b\Gܽ����?&x�4�|v�C&�oV�W��Xw��
��	�y ����'Y��tz�$�2=`n��I�P�����9�*J�y����_�f�/�N�n%9KJh'������w�{���X�ί����K_f�Mk�fK ���g��'�è��:3Y_�<�=g���wE��5�Ro4^�:�/���[�Q6��8K(���P��
T�� 4u������Wky;�c��|�?W�\��~ν��q���j+2������J_�<�[��k�5B4~$����ß���Fa/�gg�k��W.�;vf��Wg%�7��!�rh#z�ש�4�ͻ#E�=����v���+R��B�w`r~�`