XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`�Ү[w�<B�Q���� �2B	# z ��f�gp��<Pz|4"2���{�0ۡBe�k�'"�F-&�<����]�;֣j�&���'Qg�\�xf����8C WE�T�2�����W��O�o�U�"�N�@��C���_�Ԝm�����9h�Η��2=1��;n� �P���.Zk?%@���U�A��i,!�m����6�)'<?(�|���g6�ǉ&1	�=>�����2����+��څo�5�(H���숮���B�gZV4!�C\՟�߿�Q�`:����u�2D��(��)v�$��tg�7��"��7�㮐�W=��~�|6�F_�?A��xm���
�s� hRN�m��O �+k��)M�E�ɹ��s�39��_.	�8�);,���ȿH��Zc�L�=)�ߕ�Lꮁ�l�/<Oa�NMV0�AnfpW����-�n���:[딸d�X�V;]����^$�Ѷ��N���C�T��T9`�����_�g�E��^�3g4P� ��Ӛ���ՐJ�/c��A��'�V����YV @@��延��
�o�j��	���:c�Q:����%�?��7�C�T�ZƧ)ݗ׼^wc}]4�W�F��o�.��p�i`���Kץ���}�r	8��1)�?�0��T]?X-�U�b���_J1j��f KF��]eV�����&�/��`��T�m�To�����]9��D\���_�b�<��H�����G�Y�ȳ�BS���QXlxVHYEB    3dee     a605�F������̂+�F���/S�ba\�^�q� ��'�����5c)iQ�^t�?����V�}: ��"�)��z�<u�n�enȴ���-�.���z�Z�eG�Vi$%�,ŝю���bɤ�6'��� ���0V}������7��+`��9�/�K[�w�;��.��հ�Y�/�/��7؟��Z*So)J���R�&sAW��f����
Dqdp�{�6)[A+�g�9ps��#�����K�@6�QtNЌ0��[]���{��g�!��G��7fg�'���Yx������ӽ�lfJ� اDtu��(��ڛnAG��LÚ�kaS�N�~t.�ʼ�ç�S��2w�����3��vR\n}c�9`h�(D�RH8	�{<ru��..@ӳ24��'"qq��Zr_�P|�J*���9�k��ׁ��s��c�q_���A��K2x]�ü
���z7��*`5�_�`�}�~����"5�B���
6?pzW���R5o����j�H,�zۅ�[�^����ۜ$93^r@����Ar������>����텕�(69�TK�a�=�ĬE��px�'�a�T��x�d�Vw�&����
=|�92���OOOHe{D&�.�ٵD����_�zG�g]}~��.��{�z�i��;����(���2����)�o�� 
ќ�$�����+m�g��|���WK)�Az���6���oH:
^kK/^�mq45�?5��$kj�/�a�i����-ʒ���y����/CB FaH�������>H�*i�ju�e�Z+��� s�rx�3��r�3�8�&놱�s~�'���D����V��D�ښ��t�hWu+�?�(~�Z����h��}�n�s�e�'Cm9V����0�������|�O��0�^�+�r�bA�H1��'��i�S���R��r[�{�A�����[�Ӣ�@挅��w�^��,����X��+Op6���O��=<q�mωc�
�a�����V�����LV"*~�)o��\�g⑭T�=�����}1�%I���X�e�̧)h�a׼��s���js52���/Dv���C�e8z5J��<�V��n��{��X�&i&�Y�?MY�cc��Y��v�E��Բ$�n�����O*<�n��Oc�~��D�\���Tg3���EJ������u��Yhp7�n��p�x��ϰ\���,���_7��Ak�b3:�]lQw�b�1W���4�5Z�3
���t�E�y���ΩJ�j�EE^� t'u����#��@d$���Jٻ�b�WT��|�4�����d
��zl0�;`O+dU'�S�/
��|���(��Z�Q˖`\�x��X����;��A�6A���9P������<	 P-��	fĦ:[�t�6`���,��QB����[B�bU2J�`�o�ǆ�B��$���r�����o*Ѵ�'D��fnz��I�`	�}�*]�M�em��ɬv���9+ʷ��,�DÂ�*�+���T�Y���r>��������ep�]&㮗�� `t�Rs�H�)�v�w�(�%=��+:����$B�P��vUW�(���ĘU���r�yY�*4g3ך�PQi�'r胮\*N�9b��!G�x��a���-�����c�����?�SFЖ��/a.���w��CG'������q8nag8"��7��h�T~���Q�z��ZB������������T�WaL5Ȫ���1*���8�)ӿ���	;ؗDK��-)�L�*Do�]f���Տ"ݱ�h������vo�}n��2٣קC+��c��k
/X�=g�w̡�P��UÖ=սk��dhJ^��Hˑ܌T������r�#�x������o�[�P=����h2��w��弯[�g;��.��拪��`�M�W��%ZSt`��ĭ9T���O��O2�</�q�k����`s�p�����u�/���uT�38+p:83��L
j�����V����u��j?����Ǖ�����!˃���p4�{��DڦW��X�ב�<�<�&^=a�!�#������&?�-�-�=먶�>��q{���K�I�N;�	�a���[{� �`�P��KK�P�vXG:C
giI5q��2p|N���X�x�l�Ji�Nr��nHԯ��8sIjט��uy�t(
:�Ug�_a�}���͂B��<YR�}O��M�R�B�e�|��W�QWFgL�s0=�0��NUp�4$��O�����U�B�qLF��N�+iN}��_;0���Xg2�n�<�?>v�@���g&��L��6�91L�'��LJ��^���f����D�<<V���w��b'�d�%���"�I��1Wa������'�*�S *5d�% n0$����i�[��2)D&@ps��;��Ә�+��&�+��1����f�Cw,��Al��%�1;[�Ž��R��`
��{�Új@rw�-+���c�h��D���&��D�2MF/�8¯//����̽��̥��FCM�"��y����e_+ ����� �nE<�J܇�Bɬ>OG�h�zb���2Pm,2�D��Ɇ��6����CH�gn�ی?̨���G