XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���J�A�j��X^|�b��S�bB�JŢ'�1�h��j�Ќ]��e)����q���r�|�^`����[�r?�ڵ�{�̑���B���-�6�W�����R)����g���O-��3ډ�0��|���Ï;�È���V�׮I��� �<t�+�r`��3�;�\\�����Sqn��iU�tʟ@��j��L�snf'�;�>3���V��B�~��� ����9�6�~�^
�:j� ��i�<7��F�YB����ѝ�JAm2���(� �h�/î8_�z+ؙ�"YwuÉ�q.d����b;$&����"A�i1`��]��mw��������r�F�-[���Bx���'E�߷/q��#G�Hw�u����I� �vK�sиK�����7��
�*�?�`���h�H��G�"wa�A���B��HHV:��%<,F���bK�OO���:]��ĨK���_,Q�S?���'���@5e;ܻ��,1��ce��u[+���>L��d�Wdpr��k��R�/����ք%�Ir�z+�I�e�ʎ�9��25���ok6q� ��p��|�v$\y�:;j筓�
��^�=��r��z�)���;�f*��2���5L3���}a�M i�Q�Cs����)�YKj-�ڜU�܊��������~�p�uH���W$(�m����N0���[d��J�3�P;�����v��
��/����P
�G^�O��޵q�XlxVHYEB    1343     730n�&jz��ς
'�H�$U��D���
�N����	U#(�MR�������t���^E>F��3W0k/��V���.J�D�T, �c���\�{1Px�T.�q+�	��\$�0,�DL3|��0��V��{�\�값B�VU�7t�`M�^_�|;Q�&����
5�ecF��_���p��%�2 ase6�#y6i�ƫ̬h�����gp��jAz;�!t������E&��	�o�f�$��;ѩ�E�����uǨcf���ɘ�t�2��T���&0WȂ"ܽ��"�uAM��Q���8G���AT(��Q]L��|:�/աN������b��7*rxޣc�/N��׃} mZ�Gt��|;LT]3�_�b��}Xz�8x)��9m�����}���ކk��AAa�n¹Ia}�^�}
ɒ+wQl%�d��yC��'qۖ(�����:jys'��tF�Hg�,b+���@�1� �Y�~�΂>_�EZʮI��?�?nx���Q%�A0 �ݎބn2�V�;lc��l �̮6Mz�M��-�j����@�����?ȡ��O0eC���	��e���T������p��gx�>�}��(Oռ�nr��?�v	:Gq��i0�/t��X�T�[w.x�y݈ #�+��b7�9�o�����7�\�}71�W����dø�|�|I�ʙ�hr��G� �]=��ou�J����2�SEK��ZK8��kP��J�Z�����D�U�_��!�I��قF�1�O\���^���x���Fk�_4F�֑�C&i�8x1��WE���~��������_�D����=ީV�)Y/>������.��o�����Ծ���#��c9"̿7�F>��|��pBeZ�?��L�O�_|��r0�rG)��!no���f,�/Wfa���eh�łN��_�:^�&��/������6|�G�3�����-ڂ����p��c��t�G/K��AY:+�)ͭٗ�D��Y�y�,�{p�5�*`Qϐ���eH	��۹9�iO��)ӱp�2��xY�h��N��i���ņO����e�`�v��v�Y{�u�Er-е���rc3�q���+�p/1���}�uL�+ �~⎤~�4Zpe'׃��b'>�/(_�:�!�_zX�X�C,ƻ4��������n/l����f�T�d+:H�9� kps�tۚI{9���HU����{����zQ�Rۙ��&&?�׻�+{�n}Ʈ�k<^�m���r���� A�̲wX���usl�s523�N�JclBj$p��f��y���9\��f�P�?.A87B\<|>����΅�^��R��4򿤴cs�B��doܚ�R�ΝT� K*�C�D�S�Ww�&w�e��^��;bؓ�H�n���ʾ[�R����3~�\(���?�}�Q*ʸ�c�jT�f[J�g Ƒ8I�$�*?juE��.LZ~T(=a�&�5�G��Z����D��T�EŶr�,Ss����[�)�
���;��l	f2v��L���0�0pA��Q9h{V�x3�#��52�4��YY��F8'�1DVg�*(ձH�!�3��E�c�5$��Q���r26HI3Ğ��)����G����ia/E���7P����F��;���6!��1���Ќ�>�X�CYTV�ĝ�5�����e�\���v*Ȭ�D���J��m	*�PEysaزgx����Q0Ԅ�%�q�z�XJ�'f������'�{�ýS�K/�`�1GI]:7Z3,��Ŗ3vRuK�,�b�O��5�-)����Z��P�WJI�bYxb�