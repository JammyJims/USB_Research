XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|)oe��ʛ���T��5�4^��'��&�-w��e� (z����>��3�հb��nl�6����j�Ĩ�.j��'�K�T�n�x4�I��·��ۑ�jc�0��K�3u��`��������(��Sn�0�{җ�Π��Z��O�LB��>�����I߽[���UB�(��>�,�5h"w�b����%8Q �A*�Ù"�Kz����?��[�EZ�+���<�@��[7T^|f���*<:�u��q�H�D:I]|��>-��AV|���z��N�_�3���fXav��l���P�c<7�a&��c�p,�R���^�.�y��Ī ����� �����q��U��D>_a�����Q�EYbє�� IF�RR�=��v�KD�@����M�G�~э��7ở�#�䩞�P��k��Pԙf�&�X�o�]H+q,�\H��b��#�����|��;]|�2L�K�fJ7.8��D̷��	���_�v��CgNMԐ&+�5���N����B��c4tR~�Vܲ�������os ��'��9��+F �JY/x���6�\e,��D���抔X��o��#�cWzBO�E�#��IFZB�3�a��%��S ����6OB&��PP1B}�Voo"˜w�u%���>^�� DffD{������9��e�(Rդ6�l<�}���x��"=݄�6�i�vؙC�9E5&ٗs\W'���1̪����x"��!l$<��?JXlxVHYEB    1b52     a10u	(�1Bs@Y�4a2���F�{�s�k�'�8o�9����k���������
��C��*���s�ַl��ik:�k	�(���z�:�yv��b��$�����~�|���E�#�=�͞�7�D`���t�|q!ZR��ք<�����=��0��U��m�f7��W���Я&Ø���=<�| �=`��c��Z{Rx���NW)� ��������]�֘�KS�q!Cs��bЖ�B��[��
G���x�6J#�o6��u��J�l�z��W7���@Ƅ�:L���QXg�%u��eA�I�����e�1��p��%�;����]�z|ѓ�~�����h�ԣ�}�q���ި̝\�c^�f�B�dȮh��axJ�e����X(ku��6�qj*����5>�֒2AC'%�.G՛���+�?����9Gq�!)��w��(xc"�'� C��LG��w6N�ڌϯ������s��+$xGw��:$�I�#��Z:喙�Lᐢ.�w�L\n �P��P`j�5���R�VܹG\�G�iOK@�9�7 c��@��6~�=�+sM{7���Ë5}��\�Z˛�WK$���v��Yg���ӒD�g1�/��V�w{�������(3�}�d��	昴ϛ�O�|w�+����E�3WIr�
B8[?ID���1�|�C7��
x1S�G�N�����?��ʭ"^o�QJ��i�B[�{��9�S8�o-�Q6=�^��CMI�IP�bmИkے
�*-yv+kآY�M�3��|�(���FA&�K5��+����kJ�!�Nj���39�x�B�@07�K�lI���IUl�ҳ��!ӔG�owHD���]�J��f�!�N�sR��!�K��_W���]�y�ԟh�j��1���N���# ��sd��,����S���c�6���~�V%s������^�c�N����DN�2ʍ� �E䰉��o�'���KT��ͫ�p�P�mӔ��<�-ކm��iU5���i�1ܑ�÷����G��v8�],�ƪtW��l�q^����5-'4��jB��}p��\y�C	[�t� �M��#c%O�ײ�����@��Y-������6y�^�~GW�bI��54�m�����K��#��ǳ3����S�p!]t�r��?Y<ڇ񗈎_�ǃ�~�"���5.�`���~�C�d��ˏ����x�Wb�����r�j�L�s�E���c�����+Ԝ�������7�]4��e��0��K�6Nk��h���$K�e ��u�-h�C����z��]�)�9k�z�}T�B��rc�A[m�e�8��'��K�7֍�����YU@��1��Ɠ��#��ܿ�E�1�g��Jx�:��U8�'N�eF-�v�B3j�&�̊~d��K�|�Kq�/c�Q'P�7�ju2M�xQ+�|���֝'�����̡�v?��c�nr<��z�>4�te ��p��Fút��C�a>Do�fZ���Ĺ_)F��SHG�̛�|�f��M% �anו��cYj�0y�d�8_�"�@��I�=ۄ7����0Ó��<�i�ҟ$�͵��Tikx�W�f�� ��/���d`j���_v��X{@\�eF�T��]�]�5H!'��,J8������o�;#�I:0���vׂ�{�8��AM�T���=N�
s=}�g��FF$�쫶Z�a��yD�7(�����p�� DY�a�~�pЬ��|i�Ѵ�.�%���a�u@�0p��l+�r�۹T��t�Ϋ򌿪?:TP..m"{$�|���������1��M�ZNdV�e��7�!T��ЫȐI���˫���.���BTU��3+�y���H��*�)���nir�/p�,wlt���͌U��~��#-W�ȒJ �@��!�c��+�b�����(ERY��0[ pw{�&��Y��)d#�C�M�n�;�q��R��Y�IP)݀���3z�����P�f��U�K�{������,�P�Ê'�t�fER�hj?�����~;ecF����Ki@;����+��T2��;����c�~�a\h=O�Koq��K K�Ar!���,%�M�E���% ��[�B�x��J.$��b򄚶:��F��<a���D3K�7��u\M��úNi�|Dy��U�9��5>�f��mӓ7Pܠ>;Yg��/�=�N���d���r'V��,@��e)����q��L�&t$
���Zw���b�A5��{��#O��+�⍱�\�_S).U��R���yx���/�)��fx�n������D�w:I@�&ҵis��{��Q�l��h�5�f~�Lc �*xC�\l��S�W0�"I�7W4�,�ۄ�XԺ[�4u�q h7v�W���N�L�#�}��Q�.UY�r�U�_�G]���H��rpJ�c,�3<��j��>�sAw5� �W�W��-:Zգ�.c��b{y<�����Әq֛.��|�3Z�j�C��7j��Bs���,��B�h�[�QЃpJ���FR(��po!�|�O��ݬ۾�6V�N� =t�aSB�����)���