XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	h&z���,mN5R�e��Qt�b._������O�?�Da�f��a�P�����-��q�W �>b^��G�J�}H �ed�LV���
!�R	������h�M;b%W�Z|�^�\φ(��ߌ.��Z-u���ڀz�	�uE��K�/��!U6�/�V����K����y�7��s)�+EX�����s�U�v�p�M�Jz��E���Vt�l��v
M���D��'�x��jKS�d�K���M�@D���t�,�.�Yg�z��*�x�eٻl�y�W�n��\-�u�BQ^Qm�٢�~>�<ȇ���v�bپ6ti{��|�̺["�+�:�<��r�0&�����:�=_H,0Yple�]�*W<5�n����h�i����wi\�7��N��d,��,�f��<�J'`=�i�?�~[P�vm��-��G��k(��x,�1�qc���.�t��u�h��ע+���8� ]��u��J����
E���й;'��GR�#��~�we嫗���c���/$�fC [�J��8�g��9ǲ@F�F�@MQ����or��Tx�}��#F��:6�E�Rͷ�䢁�(���#�SY�=�Ӹ��C�p�����-갧b6pN���ܳ�Q�ɮ�]��Њ�6�lNs\n[wJU�$y@���t�O�P��e n+v���lQY�P���i��X���g}�wt��lC�:`����1R�vտ�a�=�0�=[�ϖ*\F���5���-�M�a�����S�U��j�XlxVHYEB    36ea     eb0a��9�*UQ>��f̻<i¤坒�\��OA�Q���-� �W�t�G<��4�1:0c/�'�>2�l�������ݽ����oAp�U�/k�Ƙ؁Sג���!s�
R��c�2Sm�dH��|4��I�~:���9����lm#���*_ ��>��~)*yb���+*h�Е�$qW��m���S~k(U�6m'����?�.{h�2A? ��e�I�  ��\d�e	�S�B�E-�m�Z������X��*�s��X�	7�-��Ak���[� �r�h�ͩ���C,��o��-�T�1R��O'3���M��ej�[�:�6B�諾����_J5���`nXd��DO
<
�K� �*�F^~6�pܕ���cxr�`�L1�`�O�.p]��_����٢rЯ��6p X/�z��7�W��J?UY�Yl���M� �.A�S2EÅk�O�2��ep~gd�d�,�7����H�%�P�������X��`�*-�D��S����*/�X��LW�h��0"�\C�����C7���0���������+j};F��o�cJ��f�.@�X�SY��0b'V���B�>ǈ��Å��4���fP���9��6A��������uS5X6%��{Es��X��o���� IN�{��Bn\�K�_S����!�G��5�f�i�u�>4�\ۣ�trq�ǖm���Yg����o,Y���5��γ��nG�=?F��-�	ny`�-(���0�k�#������N�Շ��D��bn�ru��ڿ�$�2uD����H�� 5�d�?JC���ߐ����a]����%EX����'E�\��a�����s�����S5�C� ���;T�sm����Z'w<l�T�?�s�5�i3���=0�L��~v}hE��~�����u@�R3U2�H�?�ͲTviW�RlbnC��p��d.;�D��Qf��SǇ�kyI�xJ�%q�7����pl�^A;����9��KQ ==���7yh��ڰH8ݡէF��!'�����ֹgMqu!9(��!9 {�T��G�:����ϖ�~�{wY�6�:n�j�`
��3�P����VHaD�U^f?2V����{;# �}��;�u(Y��֦K*��K���0^�Agl�|V6d�YG���5p�tF�{A �;<Il^��R�sW�F�.�-�E�\nX:��~���y�aΈ�)�Zz��?`g���`�9� n�G��K��-��F���I2�v���c*#	d0!����ʹmA�� cF�v��f��2}����`�i�'x/J��U�(L?f�:w!��_R3���.p$1��vt���|L��,�@de�2��/��i���8lG�;N���m�M��;�vF���0�4�k�����m]��XƬ{��u�"W.�7�/]A��F_��[CW�8jdqa*��F A�Pn�{9� �G%|�w0��
ZĮS���+s�G�k��~�y������z�A��X�_&�cd�p�t4�
(:V��Q�����M��\q�$�n�2�6P��.Σ ����=�l,K%�p\�y WJ�?3*`z�V��O��4yD�n�c�{ �'��>3�r��BKQ�1��J�&![�r�h����4�čI�R�Je\����
P���&�о抍q���-w^4A���s��q�o�h����Э�.-�I����k�k� �����)�#,��>z�[R� /+p1�!�<���nVܗ���X^ԁ|I���ziQ&�'��"���ӦdyPN�M�G�*�t�Iy�����%�(��C��Ї�H�j��%��K�E�2oF�A
F�Ȣ���*;�q1��D�4[�#[Q�3g�O��Q�~��Q�e�8 �Ht=�Ȃ�-^�p4�X�D�I�C���� ���b��"r'\�G�EG�Gw�/��{��+��W��<jy��&��j"=�^�Rm~���<���6���g�����F�J"9������,��g[��G����4ح̜�{vt������-e�:'m��f��$�g��(��>KAv%@=K��m'�h� 8��Ү̶��IA���>L��a���<�y�:�9�rWxx�h�)^����-��|� �u�c��	�`�'��tWB��*3�����(t�O��E[�ň�֊�6|�y�Qkg�����x����c?��,'�,�ԄY9�Ÿ@R�uI�w�	�O�YYFJ��k��؊��c��/�"��Y)I}ؠ���F*SV�f�ۜ0P�?g�M��y�������<�W�"������������ ���+�:���:�G��W�/��,�Q�����X��R,M�ө��)���>��I�=�iz1���y/J������U��W�������*�7����n(2�g:������a��h~7�c���Q+�O8^Z�<5��,����!�D% ��𾜍_ҷ�{�N-�N(6b��t44I��fb���05;�BU�6�:b�J&	f�`�bS�����<�+�?�K�ݸ����
��n(�F���N`���&�F�
Лz"�(l�p����6�'w����h{xZZq�F�����Mq��]�\���]������i��8�nr
n�'��.�=��CKHv�~O$�廙��F����iD'��hG����z������b��n��U�؆2�(Ӈ&� ]z�9��	c�n�$��R�X� z�<�!v�}�6����&H��]��Գ5"�R�����G�d\���J,#η�~�[Q=�M>:�̙b������6l���k��!>Ƃj�܁|9iN���; E������{�^~/�]��+����w?���9W��s�o����b��8�S�C��r#��,�q��\>澂YMέЖt����_T��X��*��I��ǕV�����V�gT�����j�G��&߰ť�`V�k��HNM<-QE\C	���79�����V>���x��Ͽ�����$�'� =�̉��~k/\s��ka7�]�ُ�;�&6�V��U�{t�*��'_���Hӫ;+q<}!��&�Qil��T��Ĵ����ȇ��zѥv�� ޾�-��t�P�Ȗ8��e�L��6��j�\�T��L�@����t��ӛ�O�sZÃ�.E��X�w�QƼ�v��3J�.9�`��ar#��̉�p��;$�f�|��'4EF`�ֵF/^�KM�����LvzZ'r�]f_z��54s?�z�~��UC��߰�p�[�:���/��!W���[�'b��p�:G)8m�d�,�ISܾ-x�|��{���4Q��ʲ��'3�3�X���u����Oؽ?�X��Q�F�{��#�~��h� ��}�s�Gӊ��䔶l�u��`�mliC�cT�{��؉�i��6|˭���c�a�M�;�ƃM�vG۶�rM���I�����q��_��������L���8���+Y��xû���A�+#�����
c�.k���Wͫ+�yci�� d8u\�A�c'�~!�j�3g��7\���[N.�r�5I�wx�u*��c�a����{`��@�R��9e5v�]�R�����>خ�8�A�±Q^('D����/Z�~�"������b�����j��RYp��X`�P��kp6E�kT��9����D��`4[j����U�aR u7��:&�'-�L��:�>��>��>���k��V