XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b;�K��
~A���+�t��{��:��<lU��ɏ6��rՊ��*Pi>�ʧN]���\K���U+"��Y{1x��
d���s F�ڔ�*�5�z�n�Q�ZW���{��J��s&xB����y �����UHs�S���)��i?�=5|d,Q��v��Na��bl�U��B���D��΢�eC�	��2�E�|J|�1ب���b��d�?��m[�ӌ�)����x�Nb1�	<�h\t�RQěklZ:ZJ�({���MY���n1j�ݽ�zF52(n�G�+2�&ikB%�5��`v��Ȱ���~�i�����Jx��;#�k�(Z v�P�B6lU`p��"8�������2h���I"?�S��l����D���!��x;&&>�sW�d�<xI�n�%ʯ��#�I�n�a����b��]q�p�]Q��p�
�2����;p��Y��*7��G��"�b����k���o:�5�1 ��#��ݕ��{|�#D�@n��0T�f��Xl��,��T{�X� n���C�X�ȵ��q@��S��~� ��*�����.Z��Ø��#�$<вw&h���aU��w@�&�:�3A�bʚ쏿�a��nc�C����LU��Ѵz�@FK�c��[I���v��O��ČB��%ն�����^�L�P�>�	�HF�'pI�������"�� �y���?$me�V�ɐ� X��Pe����՚�Gvz{A
)@Z�����kh,�XlxVHYEB    1680     880X3-]�J�f�T��Q�^�������(:T/ZD�j\Z�2|�D����~���Y���]�,Ĝ��7d`6rq��N����{�[[+�R���z̑7nVB��>�D�:�njߤ�T��%���߅G�`�^����Wf�B��f���2�c����8ny��c�MF:�����uj��c�~P�w�K�,izn`B��Jz p�(���vΉ6#(V�H`:��1/��ytI �M�g����<Cĝ��g��^���7���htd+��>hA���;`���C�Z�*���(u�8gO�F�I��2戜�_�)^͒Ț,=�8�H��
F�d ��4�����t	��+� �)��q<֪��L��U���`���N�M�u��8� O��9l�6���O[{��g���A�Ú|$L�����㻧H����~�RRJ�(,�\="@����ئ��N�~�Ɓ�m�R�H�@ �4W��c|q���ڮȧ�ݿt"q��5ը�}��̚��Kary��)��([Oo�(T��,���j�}�
<�]2�G7�'2��(
��l�/Sf�"� ��]�h#^2���7��ŵNU��\�N���y8nܥxIeEա����?��_P�M\�Os��fH|��H;$�jw"Í֪�3�u����\a�� �Y��D�!M�ԩ�6�a��Ok�~IJ����?�9�D��.�Hh�t��`�Ɉ�e�
���I�=)-W��>J37��9��T�8:q��၀��x��O]ta&�U��N�Z���e�{+/L�<b�l�������k�E��Q�@�3ւ`��X�4�6 �ͻ�7���1,"yh�)S���)��G�R�!C7�D�{��]�,�'%:k]jL�ϲo�����Ċq�������Z������t�d��k�"�����TШg����63kϯ�2o�#�HB���V��2!��UTo�sC)�a-g�n.O�2�=1#@o��T`(?�L��a�Ml���|��7�kQ��8�[�V[���+�vM�K����d�w����ly��[��đ�lμ�&sE��Qj���e�?���1�\�"@j�א^ʠ���ϰ���`�_.���e=�`��n���5�%�ڂ�ƛ�[�1�N���B��W>���������G{�||Oը=Y���\��0�OA��l]��������eo��	��H3��CFn�p��IM��0��!|MU't�]J�ң4��)(�1o)���O%��*	N������J�i�'#0�Cq�-
1x�A�.�>�w؉Q���矫��bp��n�W #��)�ӽڏ!�M2g�ǂ�WsW�����M�>敨�5�b��VB'��[�B�4mzF�ђs��e����S��a#40�mZkUM�c�s �b��C9�?w�zA,"���\n�Z�-�pm}��D)����Aao�Y(�r_C@>@���CU��<�rk��,�xFi����kh��ߤ�W��9�(r�.�=s��i$~c`cxҥ�U�%)��;"�rK��"�[u�,�,7 �Eł�Џ�b�ˋr������#UqU���Qb�;�;�5*��)��T7-4��,J�=�7I����w��k��P��ϰ�GsM��[oa�Z���,e�#��:P���{S������d���u�4�����a��%�>T�x�}}��G"K�V���M�ԃ��6%r�T�/��t�@��#I��U������}m�%�eIp���5b�6�:K-���*��;�Sn�����h`��g���x��DesA�^���s��9�UN}�d����̢��+C5�rfK�Kܕ�aJ�W�8aā�2��M����˃�ԨBiA��y�"���NU�Sm���!i^p�Z�f�s��5R���?DD�74eOrzO��3��ڠ�v���{��u�l����o�����>\{w&��4t7�@B��i�%������v��9�WE��'��/$Zd�p`�;������F�2��I@N�����6'h�Gg����s<1ɟy�Y�6��L����r�:�@M���]�A]�=E	�x����lf� �����1�ކ"@j�m���`Lmr����$~b6.@��J{j