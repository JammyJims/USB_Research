XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�}�3�)�Upx~�5+98>�bG�@S��f�i	 ��k-߯@�
��vǽ�D�i��޿wq!6��=�����^j����a�73қ��"q3�U� j�:X�� t��n�G��[�͘��j�6�.��pti���?0�yq�Ӑx̺!����C2qw�����>f����T�Y��ƞ�E��vt i�D����#���n��p�D��p뻢���yu��P�d��:��S��4ѕ�)K��G��qu8����﫡��Ϟ��֤��)W�h��0�H���Rd�i!���'"]sPp�l�+b�Ңb�����m�ͮ��h�l\��fƊ�{0����p�L'�����w�[A/��=E�BS7������W=���V�F�'��+�ࡽ#�Cz�4�\%gkeɇU���\��]��~"-�����u�ē�8�.H �1��t,� �>GU��)����� K:2�xAM�yd{��9�E=L:�k����4JV<\:̥�� C�QF����b�%ѮW��m�iĬ4��
�5���c�c?��ӻ�e#5����
����Cgّ��	��xܫy N����b���$
�yjKn/�5���O=nʘZ�%�A�,Xr!��f��=�e�>�y�	�&�K�Xn�}N�`r#ĝ#�r0�%� ��dC�d�wc���]:�KG.�=Q�d[�{1��-W8��Q�\6_��X�(��;��)*��_lT�pc���W���'���W�n5i C�\XlxVHYEB    2bdd     ca0��ݚͦ�7�X�m��i��)����	�]0m
��>�w� ̙!�5��ow�*�=��"I��;>�4�V+P���2��.c�\(/�Ρ\��3bJo*�T7E��7�؝H!�������}8�T�E�:�E'F���3�P�^_�`.��*��M�&��K)]�>�z֣�L�[�]�Jݫ}��H��Ҁ���d�.F�m�9�UΏ)���(O2��b��������U�;]�f�ډ_6Z�
ޏ�%��e��b[�wj@�`^Ķ��]�K(�7�<�}�؋�~ ���f�8����#j�����Za����C�/�>_/l+����]7��9�ĝ�E�sr�b������TC~ �w�[)G� Am)�\����r����J2�b�P8��5�o�sl��R;�v�D�M�����0]���\l����������~������כ��b1!�0(��T���c��%J�%�ÑzF���l�t�[<,1߾�y�YR�a�I���nb�$Y<C��������@�e��GڰJPMQ�ŭ��&�p	;������{;Ǔ�a�L�_��P�WIN��t��+3�ΝM桇f��*�_�fL�Ph������nxD�,P�m><~֑�~1����*}��f�Sm��*BHe勤3%�l���f�Ȗֽ�,���BH'�|\$xl�	:���c���L�uy�Mg%`B��SX<W(����@,�����t���k�Q"�@R������� �R�\�n���f���X�('��2WqR�:b33KC7��ַI}OZ6 4'g1��~����c59+{��c-F�UYꙕێ�ܡ�E��
�K���N��d8�b�S%+�'0�s���)�U���2��&���W�]�K��;�%VX���_
C�ަ�?��(��^ˈ�B�9zA��T��϶�s�2^R՞-n/����S)�>m��0-���������憙xz�7�ţ�
bӕ���,=�$�6�Y��9W��！h�x8p���Ac�!�w������WW�����į�����6��
%��W8�8K!��e�����ͱ-����`���kB&��Ѓx=f��$8v��梵b��s�&��$��v�Ɏ������n����&�����gҎ��2�����=��!��4| %�g]8�؈\w���A`�S�� �n��(.<7t��|��g�Tƨ�&9['!f�,�~y�UØ��r��oޏ@�@��?�⽟gEL�����W�; ���;9�gE(ߋ��of��:M�d!���n��w�˕�RZ|1UF��T��j6��~u{��Mr�i��ఽ�����L�K��k۱\A�v�-g"�aj���Բ΃_���C�Kb��":0�j��I�d6G�`JUdj���#������E/=�{�l������t��;y;�C:��~ղ�5�p�;�*�)O���	�R���K+�x6�8��҃΀+��}�z��������/��xc�
�?���w���F�J�����Rn� ��!��A�*%qO��=��Cý��];��Sn�4jwv��-V�O__��T���6�j�R���͖j���M1KF���1$X1'A2t��0`��{��G��_�|�4�VR�"n"X���u�.i��%����U
��!�>����T�+7��`�,D�cxo@�U�.��n�������E��Eɋ}0s[P����+2����aL���
Q�<y��O/��_/?�7�P��(ZI,@�����%�b8�{->�.��<�ֻ�y_�b��fq!�g����Ys�+n�lXF�9�7������~>P/D�C� 3�:K�y�]ھV��e�+\��6��>I13�˄oxM
����8��0B
�������|��m����x��z�@iB ��\���������t� G���>I �s�})�6���ᄿ����>��^��b���r*]��9���;�^�f��]!{VA����|-"�O�tv�8i!�q���A�Y � )�x1v�X����tE�B&P��脕�h�5g�g׋�r�×9~q�k��M]���oۀ5虣��X/�Q��Tl����r��(�E���f��{F=g
�h9��C2��x���)gR��l&&���4l�M�C��H�΄��X����w����P�4�%0��� �0W<��yw��ME�N���C�$ʼS8c��]����H��m7��1����A���ͫ�
���@�S_��2X��1���-/�st�+�Y���TqIɠ
[�2k��%+<6�I!��?S��oW�|\���j&��*R�NrO5�,�/;�E����y֚!:p1}f;(pp�4T�g(~�)�����Q��G�@�If�'|��u����6pv.�����}UӬ�"��y�k���l�>���2��`4�xV��EZ�2aXh8��;[�5� ��3��I�8}ka�Yi���{�z�P�{WHɣ�}~.K�x�J�J;�Ƙh��,{ܒ��d�p��"ʧ\��0�p~� 3�I�ۯ���������'��|��4^*���#=tҠCg{�r�`�)�m���lm���!�h���Θڐ��w���iΞ�0.C/��p�{��/�HO�R�U�6A�h"&R-�����}�xR��L��1_DL��e�|ͺ��U� u'L�@$d PAQdөC��O���iZ����R{g��d~��=�`�2}|�\g� VD�H�FX,����ߐYJ�a�mǖ�X���(-�n�,Wf'L���������C�z�p�gA^�%��;A%�{�{��	��-U�)|9DcЋ� @y�	�S�.&�x�s�X��)3����o�K[d�B�v���h�D�/S�6`��s���7 ��}�̕x��&lvaIo$��������&
��3x�>�o�1
����1m6��*��Q��B��#��6���v�]@L[��(�i��4M��z�VM�qgO�����[I?�Ĝկ�Y���%��y��������q�E]#����V9�Y��eqy�$�4D�d�P~� F�ʩbM�֦[��!PJK_i5�'�T@�O6����zGx��Ƴ�p����n�	�}Sle�&����p�j3�D�^�9qצ�+�&!|'S�� Ԝ$��J|�Q�����