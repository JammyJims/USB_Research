XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@����-�{_A���Ź�Dxz+��!C�>��F)�C��-n��l�p4�0�����4E5K��(��f=%c�����h+��p�Ht �BJ�zO��3�&�?���_�nI����l2[i-��H���e̱��g�V��8�����\�5m��Tiɫ3��D��v���Xq��W���n�ȫ�>�b� �u�"�> |B 1HfҠ"�����Ke7%/��y�o�Z'h%����xF� �������C+޳T�������Ȼ��57��$����|�M��@��Fd������@��{y�ct6H�J�3o��s�+�v �zߐ�����'��\�`c�!MP�a�4�aC,wM�(��Cb���`�[_b��sK�1̷��gMm�DMG�ya=m
<qВ �f���3�\�Y=*}g�xi�W�>��jk*iV����)��o�7d���⸔�J��f>��"�&R�V�}ؗ��ء���s��z�e������2v4Ry����#'��)ՠ�9�ZG(�n@B���*���s-|��g��9� p"B��C^����쨪�P��Vt\�,���q9�ҡ��Ӑ�^�X�33o�K҆�%֐���Fs�*���{���éϞ�E;���C�{�ß��0kH�M���8v
'ʲ���>�Z�ȑSܰoaN�6iaK=[V��Ԏι>�JG���\���=���m����(�J4Jo%��Kz�(�]K��G1c�� ﭅х|�5��XlxVHYEB    1594     8b0�=���X~:#1�r��Z���|��H��y!N���׃lJ����;1R�vf���S�f��H}B����J�,�"�Ǎ5�Ҧ���z|�HI+x&�nF.Jr�a�������s��y�9~�N��m��dS��x#��tI��F�Lˏ�t�`
چ8X�뵕��$b��Yf��t�,T��S_�fu�Pޥ��G�B��p ��U�����?��V�����_�/�4�|#hg ��׃�Mx����QZ%��#��) ӂ+�MvO��r��2)b1��[�C�/x�D�y3랻y�zO`N����H���z�Ή���n���ֆ4ޒd��eʊwt-������*�%�V����W-�Rm�$zn?���Iũlo9�p���Dq�:%	��+f�ԝ�N(�ƨ��Z�pѫ�M^?@����>���t�����I����`�nN:�+�o���E�J���7�<'<:j<�	7toY4H�FX~��i�'��J8"��/g���k�ŢD+���)�v}��T��/P�)��n��9�c�1���.����0��Y�V����=�׮ �Բ%YO���&Xp���M/�����[+�:����F}�%����S��W��z��÷gT&Ol�ӷ��N���5����8R�p���6;l6���Q.�uN`���:s�L��p�ʮk ���mA�_��,�ϴ�j�>���R!2D9�ks�zNW��@@TqJl�N�}�"I��p"Z���_y2*;EvQنc��f���m�����(��Q�{�����F��#�ꋌ>3/f:��x}�L��Ӽ��4��FY���n�5�f��vA�>��W۱	a�9���|v�&��*C��o{k�g~���~.4�����u�m�
��|�z�-zz�rӢ��KH��i�Õډt�����c��M[
 0����k���e�����7^���ٹB�������[��~�����o���n�)yғ�H�\x�!�cw�7��@��_�c9�Y��IR$@���1?ZD���:8��P�'2�ē"��'�i��_��t���R �h�1�I��P��OS� |:�:aM���bF�t��\]�>b#I"ןa�y|�:~ߜ�l�fB!����QI���'I0U�3�D�=@U�n�>���@�;�V��]'q��+�S��u錶j��aI�1s��:��	K��TS�!#��I����R��!$��Y5�j�`�ͳV�3�&�
5�D��5u��թ�1�.�k��i`Mc�.��C*Z��cW�(zo�˂N͐�������U���kL� ̱��Z�����up��i������jTB��N�#/
Yl��ލ���]��1J�4�V ' S�����0(�����2�̮�xi��j�7�����="��&O����{�<C?a��,�h4�g�Sθ#��Rj5+p];�Y�}�����<eU�(���o�{GZf;k �]��3�q��5�Y���3�7~̓��§|6q�̀.�\,ß�6_a�ֹ�&�S��N> ��^��,��P[�7k2��f���C������>J0�nv�fa��a��{px�����_�A��#����,�����u��p��j[�| !c�����^Kv�%�I��fӏ�[>����p�,�snC��.Ψyd�,�D��uҤI�2��j��/b������y����Ke�D��p�C�,>J)�̏���.��xa��+Ɏ��X~PW���)����}G#j�p���X�8m�H��}x|.Z���۩ɡ�`�����vI|J����=?�sy9 ?��h��G���)h������1��@'�0s�ܯ"����0ęa��BW��Kr�
M�b���k�/?��C�F��E��U䴃�|hRE�hU����!��|�b{"������e���@��2w�R�'vV�� �U��"���U5���m��(��y�!�~�.�A��5��iA��O_�4�w܃|@xС��g�����p�L�;d�;���q�EFg�k�9C�Re�%��9��lه{�G�7`e����C�f�_<� ��?ل�޽5�p�,�J�b�ǆ����(�7Ko�k�WB,�Fs>��ɮ����M���D�ds�!���V�LBs7%*�u��@�Ez
�s����qC�lt�g:y�j�xC��OXΥ