XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���uG�)��=T��
	���N��&Ɇd�ȡ'?����fS%Q!�-�$�� HH��J[�����'�mLG�̳�k}sX�&�S��W�x��ĞX���J��S�S���vR���J{|_���d�����BhQk	�y@�
X��l%E�sě��(�
�s)���)!6�Q\X�a��^����*>{E���!WxD)��4���o��l!�&�� ck�y4j7L0oR�mϟ��G��׫w���̹@�� ����JD�m'j.T(�n-�Ms�D�������bkk&���G�h���������O��kD(�eofe�����Z�k���}����s�i�qR�����
U�#=��r�B��s�UϩǑB��c����X��h�� ��;��Խ}9���5�Q���#����1�S����d�p�gPOkW
a�$v0E����,�C>�w%��@�fPM ^[��j�(��X��BN� 5�ЙA��`~�Х!��e�d��eE?0�����$bѪpx�!�{+*�����A��������5o�ȼQ�>@��e�Kgۃ�,���L��Ťz<	��z-������/v߄:�y��V�<��b~�U��g�!Sת�$�rD6�H>�.������TU��^[`�u3s��1]���*U���Bo^���2m\q�b_���w�ň}��UWn��O�ɬAz�j���#��}�v."�mu�Z3���Z!�z�Ȼ%e\>F�֒��2���n���񪛴�#/$XlxVHYEB    10e9     6c0�n�}������'7"p�� MZ���=���Zm�	�ϼQ���- ��I7zqU���>cUNm�dU%����5�c�g�+��&ۄ=�	+L�O���)��N.�좜F�3�!��DA�ĩӬ�ꈿk�fͩP�3���hc�(�BEO�F�z�x�"��4�_�Y��OD
��y)7�v�F��$̘��y�j��F���^�/8��.�m6�����`��JhC�+��8�����̩�=Q[�9'oX���j�쇕`�(��
,�K3���nE�Z�zt�������2
���23J�Y�%x�R�Aai�=�_�V#'��.�葉��) \y��D4����JIS�b��;{9����N�"GG>#��t�RA���!r��o�$#̝���C�`=�6��運n�h*cΝ��G�p�7���@����(V7�m�gE�r��u�!r�7$2hJ׎Pg����+8�$7w=�潄�|`G"�b�=/
�~�gPg[zw���ZV��l6�axbC0݇�"���gɫ�)]&0�ak�DK� �����tC||���4��T~	��B�s�ɑ��!��h�u�f�6���"�>��ϔ$Xf'�Ӄ~k�qy<S�� j�H�����ٶbC���hJ���k}��>uX��r��(��H=R@�sJ��z�G�^�z��N[ ���K���l�(a��M��<C9,"���#��Ac�e�L����{�f��@�5��m/,ֻ�S�L��e���9ͩw�����;>o��UY&]\�׊�ӻ`9H������E<�w�{֑3�Tp�F��N��L�"����|����0vP��o�^H���|f�> b�Ex�r&��.�+���!�J�H��^�KF%f'��}U���C..H��&��RP��۰*��=��ˋ\Х&ᓛ�TƁ���C|f��%�tmݭP�k�V&���_��*�!1wn*�ܸ]S��������#�)/]W3����p�mƯA�u���%�ʚ��� �\ .,�����e�i�y6n�&�l�DV�8�^�C��D�h�B�&F^S����P"�b�!.��B2ڐ���o�Cq9N3Bҭ��Ei�?Yն�^��-�x� ��|�=��3���J���l���,Lɇ��<po�w��S��Ags��}3q�t��,[Ş��5RTe ���J�oӮ��!�%�=q�X*�(���(��h��ɂa���o�z)�Wj<��.�Luバ�H9^��Q��TBH��f��	��d��:�W�<b����e��##&���¥cUg�0�#�Oo`��e�{�c��@��_�~ј�ڍxF���f��z�M���2s�uԠV���:����jmv~v���j��?�d8�ͅi��i���R�N��89�w�p$X�h��������P.��#���oE�	�#n;sU��)��t�i�d�9�By6:p�'?�ӅO�'Wu�J;>s���H�|�k�|$[�,`/'���E�ЊڱN+��ވ�������tTw�(G.�Xw��c*o1�!�ZO�Om5 ���#]��:A}�Dd�4��ҷy?*���;��c�%GJ�������6�I�f}�*(gs�� F�Otg0W�_ʌbҹJ��0��+�=U���$��n��t�r0��rdo19u���[���C�Ʃ -�D��(��Y�϶dv}{