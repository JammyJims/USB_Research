XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��̂�h�.� �Mp��cM�m�c��	��n�����_�Ɗq�������K`�*�^��ϗ����R#��O�
��x�Z~�kE�D�8V�ϮG�y)~�*�eͿ�������R���܋��u͎�!�,�3� ��B���#L|����x��g��dc���hAh�n�=�T$>vk���ȟp��S}�Zm���{4�-b�[��A�X�dn�Ӿ���6��r��=ױ�0�X啰,�lo������wY�G~)��d�����FX>�	b��U�Z<�vF�Fz��hu5`�n����6:�̦�?뱅yפ����!+x�Lv`$Y1:.����Ǜ����Z��yg�.���h� �'.�K�\u��,[�sb�6�Y[*i��EG�=0B��$ٷ�����B`�"��\��"��G�[!�E��Q��G���ٙxW7���e�l�<R(
�����*�\5*HU���n^�e]<��0rv���&`ޓ�e�<'�Y�	wh0�Q+?�$"��t�II2���-Ա)E��Kx	&�=���ĚX��b�*���l]_��tX,ޖ�w�!y��Ow��7��q����(o��=ìf��5պ�g��O��]�zx1��b�c�ϊn{:,?�`�|U�.���kpM�9�m2B<�T6��ް�?��{8���P��LqO�=\	�o�Ѥ}Dc�1���b-���&�k����ɦ�Sёj�Sl<׼�q �E��=�����]���P���^F|�U-�I�iWXlxVHYEB    176d     960\ˋЈHL�Q���&(��:~ě�WՆ�c��q�X#�&�������%Mz�*��gk��ڻ��H��� ���Ϯ���!!���r{Fk��c�� �md��9�>�����[��H��c�]�Y��,��)��p��G8���q��"��[L���J`ـ#�^Փ��6�7%Z�"j�4���*�`]7�|'j�Se5'�)F��ves�;��<!dm>uܙ�ѣ�bx��6�@7����S��������T���#��f�7���r���p��HNֲ�
�X^"����W�OV�6�{1&EH}����$�*~����)�g�p�?�:͇�ܩZ��(��%ݪ��,��9{3tkc>61ZD����VmeY#�2q_	f�`R��N�{����j�-�K��S�`ExH�)1��T�x�Ŗ.����ع%�{��VD��u�� 2��F^����I={���&��IzA�P�/#HwX�H.�{��
;�@�� u�� x�H�k�v^wiJ�Q4��������X��Z�����"�sVᯨW��z�c�j�|��h[W�����N��½|
vM�+���T����~*�����(h�m�_��h�݆�r�D��NR�w�=�5p��0��A
ri��~z�Y�媐~[`4�w(&����(0E�h�
����-H��I~�e�6JA\
-2]��������g��4x3�e���J��3Ҿc1�t7� ����&B!��Ⲹ~���O��TqP�2y���<p���'�f�	V��]:�.�xaF��*ō�q��Jg#�s
���B��2X�Cn��^�K[�y���7�Z �$:��W&';Q��yYA���5�ց9�6�F"C\�@=P���{u�T�x��dpM(<�a�H&t�~�k#T߄�_�5=+a}�zB���$%�є@�5|u���i�丄�fOG�ۈ�P0
�x���w����X�-W�`�x��������j��^HüV���$�tQ�g���ď�0A�Y�S�ſ�9�G�l����r���*�f����p���)H�c���7���VU��R���F���p�ZA��Y�E��A�`6�$�G �T��Ip֠팜���Ax#�L5��뙡wAi��^*��E-�\z&��OQ���:1��M��lHa56J�)uw��4�gt�S���T�]�=���.�����(/�;�s��^ ˣ�� ���0T .Z�d@���i]`-���	�9�������Xڨ*�ԯik�<6$:�&9�>Z�y�@�u�hJ{'s�I�R�;��-H>�� �����X]IY���uYc��z^RpR�n`���*����'0f}.N�4d�i�=��W2b���^.۵w�Q:�Z�Y�^`#h������~%��n���MDeRA7�����E���cl�<$�	 '��"`��ׄm���ʞ�7Hw�g�~V���JDy���ろK<��/�����(���!0X�[
5��+�\�G���~Hl�ΐLc�9[)[�Rg	\o�(�.(�E�	�{�O��=.0�|�r��H�������k�K"q�F�AQgNm�a@@��qq��,�&���&W�E~�DM�S�f�/`�_�BI��z�� ��K���������`��8f�ڮ�ʈr���h}�}e����r�}!e�Ћ�3U�2��F���^�t�\��X�����p�_S��hnD��� -����9�����h�l=Fx��ƹ�J�>	#^9$Y
0�m�L'���΃�L&�o��g|�~/�)�fY�_�߸����#Z����/,~)�o�f����&�y�fͤh�5Wɡ�Q;W!:�j(�D�S�h�/u*��J���J��fHi��]q1Pi�#M�P������CݬD�� u#�� 2܋��d���W���ц�{��8���Y��5I�Z�n/b9��>�{tΣ����KA����-�s������R���iF;���^T�����qY��|ʉ�ET���kF�]@gtA�
=�k��2���=� sDd����?~���d	O�u��1���0�@������:0��OR���ew�x� T��ٺ�>�(�2�0q�.��n哄C`g�ё\^�GA��\��Lz��N��0�^W�o��%\�C�a�B�%��¶e9"�\j�@.�j� ��/�
�I�v�$x�~f�w3������x�K�*�{��[�ۅz�!�M�4�'a�z��xT��s��������5��9�ƽ��u�W5յW�Dw���Vn�XX�Jj���jYM&9��|6"�1x��A�d��J|M[��