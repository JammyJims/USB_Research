XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v�������Z���r�O.�'('?�4��y��B��;��U�JXM���s�n��G�����	��}��`[��+��!�#�:�'�$�B���na�\�i���_|P���j�C�#��-Z����(�jT��a��NM����9����e��-�N^��Z�-�Kl���e�H�Zc�W1��*s	fmb�ɘp�@
�5IP����{#H;^�:�R�\'3��{��I#э7��f�����@���`5K�9'#z�G�Y[���=�`�7@�ː(��o�^,�4:���%,i�]���� �{�B�܂�.h�>��^Lv꣘������+�v��I[,9}�<�x�+�)"�[�#6A�˶6�bN�u��|U%�M����- �r�5Mj�{�lY'�y��Ȇ�L��F?���_s�G�͊�����d��ئÛ���G|�F���b�]k��`�U�X5&	҂��s����A&��v��-��BN��P������Ty���z/.�$����?�;�`�(8 ƬG���}���"��ئ�����kh^��^�ƕV0��G��GB�Oz>'L�߼�-���J�1�c���_'�R\�O4h��ɹj�ꌚc�_Z�H�b��(�͂�����@A�_��!ɞ�4��{��QR�-�BG�mn�[����"�¦G3 ��=��9GSr�f�}%b�x��`���TU ��:���7 ͋_�8��N��z{q�tnoS _4ь`׷ӏ�Ϭ0�^��tTh���䘬�p�r�}��p�HEXlxVHYEB    20ab     c30��L|�k�CC �AD�틹�E&xs
��CF{�N�ۨs_��#����&�̈́��߶w������'�|	�f��a$�UlfV~�P�+Ś梱ZAb��z������n�y��o�W	% ���c����NB��{.6��mɅ�<�MӺ^ZN�T_��l�$�U�!s�M���̹o�m��<a!�J��,��w@_	��=}��V�/e$��dt:�mQ&�o&D�U���.�B��sq�W��X�츤I@9����pଳ(\Q0O��s"��{��r�D=�9Ng�eva�m)m���ۿ���\�ڲ�ye7w�[��x�`��G��9$�!L���]�l�D�N��Mw*k�m������0�ƺAnFk�o����,��\����4�P�v�D3?�BT��*�g�F�k�`߄�=��	0�c
���h"fdP?3��>F���)f(d�]Sފ�`,p�E�3|��lMYP�)o@�{�D>a�����ab�[z��}Пw�Nv�Ս�S�$d��Si&�*q �f��C�%�5O`�g�J�3�bul��p?�xQϜS�B��a�bh��]a�1���Xo�=�?cD{��h�ou[�����Ѡ��o�Q"����K����Vr)���<ǟ�����]�8�u�,*��*"�D�l���� ��y�IY��	�]~��~����Y$G���x����wm��\n�W��������ۑlȟd��q������ߦG��G�pze�[zz?����Z���h�G���6��q�K&�Z#¶���+ep1�FZ@z8�3?�x���`�a_��iN��D��H�w�ve�a�O04'���=Ɲ8�����swC��j)DAU������Ւ&p%�0�\ݹ�%xL��u������~�'?'\�,��1�C��GGx7�+��d������ю*��2��I�Eeُܡ	K�������fgu����t�E�i�?�H����1Q�����;��epr����ʯy�,θ0mHJM�8��M��5J.��z���w����;W�b�	Z#�a�O����oJS0���r)FI�ߡTz�Z�FJ�}U~@j����)1��1c��$�h���%�"�}��x�� �,E�/qO>�����`���9�Μ�
a����Fz���I�N�	�b��{�}����F�q���'Y��	��d9>U[��ʂ�@k�hk���A�i��f�Ϩ�h$� ����P�}�:���?*�[�}t7Y9m�A-wb�;�T��?�����4��:4�K�},�/yfr�.���Z"�cI�A�3�fF�t3:��d1F��3��a��4ʛ2�I�N���=�:�')L��s�z5����2��6��83�v�%�
S��Ҕd�K0��ʏ3��P}A�t6,�lc���}�n����c�q(�=\��F�L��]��bS�[��}���=*���J�X���eؤ 1��Kb�Ʉ�e�*��԰������'hU��E ���a�yO=.����1���.*�!9z�sQ����$���T�z)��$
	A�:���O2X*�!Mҽf=�r�����]ȨxLg��Q}cn�s?����N��-�D�t�o��T�w���yև�h�_#�%@'V��c��	 ֣��l��1�׈���>t����$�4��1��x�\x�lv��'�}8� Ȩ���wQΟۺ�M��j���3�?�+8��3[	B\�]�^{��3B�e�h4oܫFR���!.��*�x�O�yYږ�"#���-60�Gp�d+>�0��j�kY�t���m��,?�H*�G���#�o3�]��.J�ʲ���|	*���� ����{���A[l��&�8���!���@M�\2��p���}x�p������#���T|a!��e��3[�n.����8
1���}����/�,���UM���`�.\q@ ���{6�7\7-o�60��k�ƺX��D$pCb���C�R�6�ك���ef�J�-�AD�P�d6���*B���ک����ڄ��z�å{�1�����Q'�О�;5<�,��E�����9��O/�$�@Qm���oo�|��v�V���	�&9t?��^Р]	щ���M����&�,��M�9���f;����	��� �����P�hw�mLau���$L7|���+���bv6��0H|v������d>����xf96���b��Ŧ}�����"�>�o�+�X5���ߓ���6�;��g黽 �����I�x�J����Q��o%���rrN��ȥ-��mn��,��5KRv��5�d�a���P����k��Z�HS�O����c`^�M�/<-�=�5����m����,���q�c��i�=�5`�H~�_���[+	z(����\q��&���C�!ͩ8��� vᶍ������J)V9c�Z���ӻA3�YX!�j#T)3�>b G�X/�84���˱�G���S����1��ﾭ�E�� ��!0�>SQ����va�x�YFd�$b�o���]z�������_p|���M9s}���No��aZ�GHE!�?�q9SVY�`��O�!��m�7�T-H��n?��Z'޷�5��T��]��8-.����~E�H7#ؑ���H�R6���vQC*N���1��x��>I�)����څ�3��'���l>�/����l���R��h�/��b��أw�4�Nq��$�.u�y@�G�3FRú��Q��3��,YϷ�$:��SY��T%_��(]�_b�vo���f�q#�X�w�h3hW/I���<SG�W]a^Vo��]�fO�T�#R+��I�O�{S�'!D�'Wg�h<�����Ѓ�ħ�C]�:P(����Gl�%�t����X.@�!"��^u�,�l��Iu西0��o/���yãg�j�o=�%�����ML>���F@�����mPCV��)�[�
��^�,�KsDgN��5C�ǱD�b8���(dګ�앇:���̠@���-�[��X��ѧ��pS�'�� '��OZ������ԞB��4���R/.-�l�1J&���0�ݤ�IT