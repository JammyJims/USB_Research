XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*�42x�F��?А��ڤ���[p`�z�RR���� Ӭ�݋����V*�W��̃H��EH3�/�'�����:1Q����#���G[��\�,yz98N
��ǡ��pT=���>h�̻�e��=-�[0�����%^��l�ёK��A�7KG���Д0w�2n���;�^�_L��������0�T��:`�v�6�V�Xn�,[
��da�4��RB��y��>�˿��:�K0 �dZ�pk�yWD����[T+Q'6��?E�0
{l����DN�Aql�����A�P%t��+��#�hT�zځ��?��9=�4���1�:u��)��򦒮V/���8&�v��0��q���J���N+B�D�Y��nR	?�5��O�1$>����Ҁ
�4n��`�NU2"7D��K�E�c�,�E�\�r�8��\M�׭G��uhb�
�$#���}��YLi�W�"��|�����U�3�~�,
X!��Z�f����y�OE���\�L�]ǒ���&7DS�B�KB�$.�5p���ܒ��(4䲛9 -+�i��~o�kC����e��S�l������5�$G�V�� ���H�*���"�R��!f5`h}�haG��'\����v�̕8��opڋ0Bc���et��B_m��}��<U��@}TB�j}�Z��^���4V=�h?�R2	ץ;�kdK'�&�!��2\=,�����,a�{My+M��s�o'(i^�A�̺��=��e(��=1gc��MS�YA�=�@��XlxVHYEB    1891     9c0�,{��]�
����;��T��d��Q�Y�F&u��#b����<�>d2O�Ƴ���4�绫R��W�6��_��zQ����g�`�0T�͝�>M�*�,��v��a��'��$�N���W�,�=K߾����~XOί���}/��ز>�#�	���Jq�
}GL�ˉI,*nn0h&�A�M��	Ng��5�Y��"���\�m���Fu?���4	&�9��A�e_<�ܵ8��V��/�Ч�mQ[��Ԯߣ~�S�"����l�~3ˮytDlDY���«_�Rs[�O���Z?�Q������w�� 5��M�Vы<f%9��b�8ߛ�+�2�4;����|ZE$ wyٯkg�q?�:&�ir6��)�p��ƁH��U�}:�>p�����$J��2Tb���O3�|�6�=�@��BE�	�5���e��Վ�/��ڻ�a�+��>���;�<��tiÜ�B.r(�iWI�^��Xl7p��r�K�6��A`��ǝ]��w-�L����ډ���du�H�wWH��209��p�l��d�Y*��t�@A�)<�{� 2-.�����/��V��`��{�o�$���4�k��iH@��S[w�a�:�߰w�ȟ���c�[B���A8��O6^[��0��M�F��8��Vv���?�ߢ�h����(��,⃺������Z����=VD��FE�,T�H@����P�2����K�mU(�h�rңe~���]�����Y��~f�7�q�{V�]ƴ�m�W����hM"D� "�~�"b#N$�'Ǻ>P�	}�@���f��R2s�sٖX��k@�q��-���-񈟧�߁Nd�F�	N��;c�i��e��|������������b"�n�p�G >V~�(u4�����5Va1��hS\h�f7ߟc���&�5�u�__8�n�
b����N�����;b�h��ڕW�� >8>k����-K%�Q�2��h��+oFՑ��G�TʞM^���4m��F�Lk���,7�K�����G�Q�zPݐ��(އD�=$4��:^�DqSW��:�dUc��ӻF�m`.J�8��S�_{�ښ������W\�!�?�ب�"k��#v��Q� �V3��(ܬ3�N'-P!�c�?���Z�N��Hehbȹ�G^u/�Q4��}q�)��qè�Q�r��L�)o�3Ȱ��U?��m|���\o�F]Ae�øh�@��k���?��ww�}9O,QZ�QG�o^:�%�!����Q��_(=���S�c���^-��nm�7z�X��ֿ���k���ݭ@��&��"ff��3�p�w�z�]0�Ӌ���&��V�	��+���&����fF�|�,����9| I��M�<���
��?s� �Y6�|�q�0[?�y�]��OT�!�7g��J�_�e�.3�����w�`Zi�W���0�����ĐZ�����T�|�ӂ�Vu�����ii~�;;x�J����l�|�"���X����Fe>v(���}���/���1�Uz��kpѡ1+�G-O5(d	��0���x$r�ƒ����d��`/��"��-�y�A����|f�������>�Ǵw��4Y�N��zx�ge���|.�!�_������aU��lvz�|��� ��v�Y0���?���z�#��{�@5�o�_��W��x�T�����t-S%j?��Z�Ŗ��C�;�������l2q}L��m,V�_��]�*�f�#���:ԅ'�x�` 4�ߕ?��G�8�)�3��ǌc�����<�ZCi�FDx�_��'6�xJ�x��M�nef6P�CL�]Ap;�lIx޷��Qo"���%m�BF�l:�͡��x��1,��A� p4��c���=.���ک��J�D���;j%��S�qrШ�maV����&���|�k"��ǹ��2�
Q��Ɖ��J��[���%]f�F<��П��Ŕ���J,�8��c}�L�}J4��#�n�A��Zxu��$;�d6�`g�ϲ8��Ϻ:��G�zŋ��Y�`�4Q/�@��/wh�jfҴ�gX,Mv%�3�����{��!�y^��߁C!�͝���֧��|�|��w�jay����,?Q4U2;-h[��w0C*�p�s���.� S$�v�9�TO�]�+	_���F�I#_��pY�7�G6Y�bfk#��@e���	�� T�t�0^/GBXO�%�K���K�#��yA����Bʔ��ܦ�Qy��UPf�V��f�&x��4G���P�% �k[z�*�֕W|���KU`X��5�������A�{�\��b�$�?5
��Q3�5C�s�^��m��q��&S(����%�YCK�<=uD�I�A�A���#�p\
_5��	�DQI�E��t6&�؟�U�����y��TJOyu�.Q���<3�ǲo��]2֥��1��|�D��@I���/�ω#�*s>W�Y