XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ёӡ�s�K�l�Jس�2_��҆��6�؆A4�묎5IY�����R@�B�Mд<��c�|D	A&�9�d>��S�&9sϊK�]��{Yg����!*7��Hא5$����[-���&�䓅���3KO���1�ND�$�#���}�"r)O���G@il�}=E���I!N4|��V4J�0EҞ��UD:8�r!Vd����bq������"��c7���d��o���H=�"���Nb�
���ओ
V)S��M�R䱯�ud���&x�J�2(g�:sy ��F����F�@\b�X�E��b��n��2Z7kw塝`��.���Y���O��?��l��N���w��ϛ�44ݪX�����AH��P�9� ���5,�����%�a����Zw�#T��ƺjq�|�A�W��9Ct�r�rL0�q����ѣ�������'�^�AL���_�A��@%cU�c����8���3�X���C<���@nH�6'd��>��܅Ių:7�"�������W`�����t�'~c��te��Q��P\�[�LX��IpVq��ÃH%/�f}ΐ���q���17���E��W<�6�zߦ�����\��y�������S/�pVe�t�����28�CDG(-��7	���"j��A?0�x�fA��6�'o�hp},�V��6�*�"��Pܗ}!�~�c�2�������W�����F�7����c+K����$9bϪr}�XlxVHYEB    2bbe     c70!d�5��
��`��U�L �'����� �+�f��<Vڵ�W�4m͙��c�I�
�
fo�E����,[�>��qR,��h��f��&+HL�"?L����I�g�v�Y;N��I�k5d�<��o�^ş(��.�}�2�Q��A`A�I���,�aK����wb��N�J"�Z�.�*@���U���
+&��pw��,�O������Qr�b�|j�_�3��G�~G��K֤�8�oD�68U\�Ꮫ��ڒ;2(�����I�*~���x�BѤl���q$�h��,w�]x��9��kJ>6ܽŦ��h�b`��E玲_�^�C��b}{���A�4�lN�F�c�P��Q@	��a: l}�����l��	�=�&�:��⣪m=�.l��G�y���HY��ا���ˀo��j�V�+��Vz���=��*��H�^���)����0�(�28Vi{s?�����c�F9B�"r�:IY-����o��t��N	�.��G��=D?O5} ���0�B���G<�k$�x���� �y����$��2lT��׵��N�#��|� (�1��5���,�M���,�Y#�t���K�A'�+b�`� ��<WKPAK��oۧ��M��U�d<��&/`����A׽qzˇ�X��y�8�6��#VG�%�&2�f1�9�(>�>=�g4�����RV�$����t�׷�~�]Fuf3��W�q�G*/�>�D
��	G����ȑ��<6*�2T���~̍�2���%}��_g��2ͦ�%��>[P&�|g�ѳ|O��ca��Op��TK����37��O��~��`i]�8��z���:���:��^ϧg<�Ӊ@��0>�����Y�~A��pB�a�;B'D���L�.o�d'O����{�*�����>��v�Ha��8Z�YքD���$����@ �-����u�烅8�nND���|���pms�+Sǩ�.{���p�I�����,k%Q���ƍ��[b=�ù���k.�����
wг�~R�0�Ho�J_[	�|��� ;�*/�!�z!��Ka�bZ�+HL������<-��%$���{�?#ôTh�����"��;�@��kx�9�B8Ӈ��qb��n�y����VJ�c�3g�7��]qv�}���Yk�?X�t-��PI-�IH��d��ϴb�J��������h@����q#��_�V��Fp�\Z,�V�{Q��©���Zo��1s�8>�%8��7�i���=N
Zs��d��v��0�г������v'����o��N��\�+��hDƎ����ѤC�(�r�^E�:�_���1��w��CԆqz��wh�뙐�y�\���'(�I�~�W�t%�O��6��%0� 0�#�M㫙Ѓ�R���Ŕ�,��m�B�J�N�1m��P�\#W�X�"�;g>�ǐ �"ҺU��i-3QxЁ��}m����-�l��kZ��͍/�����rb9�؈�i�������ֻ��v#rG`��
u�  4�9�r��p7h���!s۰g�kJ3�h+S�_D-��O�s�'5*�5i��u�\Z�-'��#kǷ`��������>fB;m���+yZi�.Z̤�x�ǹpwH�>�2yG��m�k��&���cvWBrw�2���_v5!Uq�p��Q
�� ��j�� �0��Z}~V����Y��ņخk�B��m�q��5�#F�0n���/�V�	��v$���F�řY� �S\`!�F�'�~yh7vZzIz���q(�F�ED�B-:��L�����9���vrs~v�ˡ��U�
w�]�0�鼼 ��'=� b}�D:��5̣g6T=`(�S�9��=9)�FfG��=����kb B\�:�qr���`(Z�_c��zJ���8���h�@4���y?}_�s
�u�O��I�O+��Nٵ��	!���Ly�|�΅3D����r~��h��,f"�ی�`{�'��=���2
C�C�'<����pZ��a㤗d�����O�͊����7�<g��8�B97S�ioL`䴩:�(�E^ƕx��uu����89g�U���)����8���8f�:	J�ρO)��iՇ�9�}�k���\�B��5��oz�K׌�Č�?��P�����"��pۡ�h�F��8}K�(��u�	�0U(���D�7���I�^P�����=�Zn�$��S���D�P嶉&p��W�!����P险�Rbl֎�ڸ�n�?�R�{R��a`�E�Cc�X�oa4� b��oJO=Zfyi�*�T2�kb��� p��q��9$O�#;i� ��:n܏������ʓ�Jǂ�ҝW�b�A�ae�$���ù��3ăE2����4��A�u���x��F��-�R��C�.����Ʃ�8�'��O��/Ո̞B��l�c��R�����K�vql��䥈���eS��ɓ��qC�+C4s�%C^j6<��"�&" �A�H'����&}� -PH� yĝ�1�	�	�r���Y���ا$M_D��A
��f+Gt�Xqн�?J��b��@Ï�H��y�)q�(%'� G����U�J�������#�o�ݧGz�wU\��Z���B��&�b���`V�)�#�bY3��S8�p�Y3���jSX�ŰTK��� lpV�;��b�ͦ������8*�Wڛ��YP�%��x�Qz�߷���v�1�8��.r2� ����<��=.�OZi)	y��	\V\��+��	��kǛi�W�	�씐Y�ȣc� b�bY���$M8�ށ�@��b�{�A�BE��ƥ״(rpX����C_����P+�a�A��Wa!>���>�@��Vh_G�P�N�8�6�9I�&Y9�����.C����Z�Z��M�`�WLf���$�_��]+����J� �Y?�^*J�H�=u�?Ka��R�(T��ɱ��"��-�]f��u����_J^W+eU���]�-4Py�}�g��K��h�� 7�Lj���|�/[�T �[�m_���f�)w���,n�Zs�<󜲨pr�$�.���	��}	�t1"��Ww�GIĦ�
�n���e�Sӗ֢�� ȡT?��N