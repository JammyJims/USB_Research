XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����j}��qX۲'+�@j��N�p�	��U��4=w��ߌ���������$@�P�t{�M�<ĩf�B�}*ݏ��w���)_�cW�	}��P�4�INno��`am����@ށ�?��@v����x�:ZN$O>5���m�ݕ�$q8p�LF�#� ����EVb[Q�5=*S���зi���GuK��4��={]�x]��iW�6���@�r�˂��b1�$�J������9���ȼ��/����'J:��tw&ZSr|�K�Ԙ�x2$�Bh҄ؕ-�s�ϺbE��Vk��w���c��ũz��x�a��?���i9����������c�[���Ă؂bDl�ʃ���,�����8p���\ӳh}���U�ŀx�Q��Ez������ȁ@7���t�!R���d@]z|�Όd�4�U�z��+ҾOs���9��:���oF����3v\��~�[#9�*������^zWu,��m4������[�l��b�@(��4&�,0��n����`%��bX��b��T���Q�@���('L��I�?�٤-�e���!�-Ѭj�p)��i#/�v�_)}>�0�2�>#7䷗�[�ۉ ������Փَ�ꡤ�`�����=��0-N;g_�1�p�HZ��Z�Hq��45��-�~l��� �N�q������7���-/�d���:���m����Zv#cm
 �w��2D�h:��s�ӆQU@9�Ck��$�����=��.{9��ےXlxVHYEB    b306    1ea0��߭����b�7֫���U�NW�3���bkA�o�|R\��"0�{K��P�)BKG����ݸ�S���	����M�He�C�ӥpm����+1KǪMdN6�����o|�rT`�sC[�pRh:w��u�މ�魼�ƞ2��Q�Zj'M����c�iϕG�r���^nrw�_J9vtg�G��D���yi=�Ɣ�ُ��X�w�Z�L�%����_1���Tn�����~?���+lH�F���rQ��i9��^�و^����� �ˌ!vcZ$�kT�{#(�����s$���d�Rv��k�C���wW�p�s���Z[������kv�3_�B��jy#I�������Z�"�"��)_Aat5�G� %Ai�&D�Fh͇J�~'ӗ�Og�~�[�Ӳ��.�$��^���5 ��ߺ�y֟d(�1��M�|
8Z/y�����i��P/�:ZB�/�
�I�����?��@\eAY��0��;{��� ���h���kF6L��D���p�?���#�\�vTo����"��9��|�?���(2G��]ږ������W}�%�_�u��7�q�'L�ڎ�ؿB��x/i����C�T
 )�װ>w���~S���)�{����^LD-�X�o�`r[��yV?5	������=���5$M-Xi_��q�P�/>eR�C���K����C�}��� !m���0�(. �ɚ>�
��k����T�B��=�n��NxO � ��29EC�<ɶ=��kvNIC���h_��:���!����'_(��}*Yt:�ɬD���1�>d�*���R�Y{�������!H
��q�
b�<�HF�R%�ng�ɧ��&������R�#�����36~����ʒNt	y�t��(V�L�D�V&�!HG:F�� tn�I.�-z��8N���
���v������di�=�]>>���~������MbC�^�l �<h�5�QQ�-�� �J�эֵWz|n�W��|�	����?0��ƅ��Ŗ.�h�s[_����[1��'�a��K�[���D�~�d܀zkC.��/s��L�����:��.�)��u����u�*|~��Qe�ɰ�b��m^/�U7Ė[��ox�E^�wo��!�<^vk�}�Gz��_�tſ*�W)�ĖWud���m�e95�es#��ɭ���#���>�!k�U�`=�6u���l��~i�Ҹ�N��^�nA���C�� �i`�!^��i�S}��:N�8M��q1E_�\�0�cYfN��_�1�Ip��n�D�t)�"��9t<��-�12!Y5��ϊFTd�yh-ym�)�Y�W���rɱ �N�"!��딞�Q#��ٶ�Y�ML�{m�D�:\%urY���g	^�FU8>i��H�0kd�t��q�M�,*AM�'K	�Y�nTa�m�4�G��=n]��{>3'8�Y �w�bɾ�&�1��\��<�{u�uh[Į>Z��,�\�@|s>I�v��R[�;I��\��ݘ�nm��g�`WT�����܈/S���"*�6C��-�M��`�=���c��܋g��s��E��<�2������� �U�(o���,5Vh\(V��f}�N��!�A�IX��[^��1�Y���h������0�% =SP�1�N�N}rk�����AY���6���Ϳ?���=�vV<4��s�)'�
�}ր��e,��u�քF�+d�;Zg Q�G�La�h"V�Bd��%��~y?����gV=@5;S�<�%�bS��a�&�/�V��5�8r�rV��=�5(h�!� _902h�!PĢk�:>�6�I]�Is�Q2GvTB�_'�H�N��:p�VQ~���z��$��z�\�s��2a!N2,t`���"�٦_,s�z�#�^�q�Αm��fҰ3p�6������ql�T�ڴ�8�]����к|x��%�A����vQTf�&n@"��T5���h�o¤�(�Ճ���o�\W�� �"4U�G����H4����zP_���D��
>
��J������F�݊)�3w����Y�?Q��8���;}.�A����@ @J�LT�)Q�����3ם�������Ū�T�$�1;��
�������33j)��u`jRb=:`��nJ-{7����679&˥��7IN�O�,���G�˘s�^4x���B}��Rr�V�\6��G��m`���͚ ��M�?�%�7Θ�{U~[��͔��9��R�"�nH�z�%������T��wA���n�u\�S���$^�k&#)�룃��M����h�6�$@џ� HuО$�g�w�x$���u�}Ed̋&�6e@@��\�yY��֭ !�w�'���JD,.�_1���#����`�V�崀܅DلN�w|�W#���K0����a��p<ñA_o���
�~���V�3��Y��lZN�pY'7Vm�=�U�����c��ݏT�R��QՎ�Q���⋧԰:��c�@�{�뵧M��o?J�GA@ٳ�Q71�Ou4���-����Sn�KMؑ�����^k8L3�Я`38�S6�Zc�o��}]<��]|��S��=�׈�B���_ZѰV�aF=G&>��چ`��q871��;/oj��߷��똕f����}�����ku�^����w�EϧC����M���z�f��(-[�C����B-R��c;���H���C��YqqG
�������:���@)���Ƚ�c�#ќ|wOHg���-�d�b+*ʒέ���투;i�(���!t֐����i���[>ܖ#�X����N}B<.�#�?�81�Ѥ��� 
��m�A��2��lʰZqh�!2{HU�
~�7���8/I��5�����]�����t4G��{<x*���R�����9��@�B��1I�v$Q.S蜕��K\6�P�3���x��9Z����U׽��Ƶy^�WѢ���nE�C�/)�`-8�;%l��v�nX
�p7˷A��&�φb�����$��U��r��I[4��o�T뿋Dhl�@C�j��tk6��z\�?M�c���r��̷�^m�h�F�f���a���5�7�֤WA���/�g��qO<i�6�wR��tO���MK�8٘&��1�W�ڠ;gѠ���������7&��dAS�庤�?4I~���+ӑ����V6�[�i���9c&Z�����LJ^��x���Э�3�s����d�n���!um"�8Z+w���Xm��?D�����[�ٺK&�5�Y���4����uu��Vt@
�o�\Q�Qpw���nO-�8	�I�#�P&u	!������NS^c��	F$L�d���^_�5tH�K��qG]m����4w��M�)�|��?� ���D��!?0PU��V��1A���(�w�-H���"V�냵���q������U$x��.S�����]e���[��c�s�LT�x���Bo�S�G������$��K�T���y	��~�Va�>�EmQ� )��&@	|YZO�����9�/W�\m�X���-x6���" �p�9��A�p�ZD��Bo��a4����f'�,��`���օۊ��	�`�Ё���=����O�g����E�Ց��#�D��}��V�:Q��"��M�7��*�d�Z���o<�ept��Gl)g��#����a�M".5��>�I���K�֑��M��*GC�k?[:��vϊ+;�K�&�v�z�D"ʴ�M-L����b��$I�H3S�:��}�V�Ͽ�VW�
��,��e���]����/&��"2͍��� P��ǃ�<yu�{��[q(���r���KU�ւU�lb��SJ�����Ƙf����V�6NGǅ�i�(�L�o?�vG�v�XO
�
&�^�tx�`�=nMI?����x	�-��,�g[�����k/#��0�8_��5r6��F�4$*��,W��+�6qI��f�A�_�ſLɏ�̒w	eeM��uo�֋gX˥���\�ԍM��Q�Dx�H�t�U4��8���������M��Ѝ�_��O�9�8�#+k�#��mLK�/0=�����i<�p9�1+�$�R�E��ѫ��k|M^y)����x�K��gTJ�&p0n!_V���쎂�3]���v%���^��h˷20�����$~��,j�}]9 0�ԃ��[�}cBgn^��_&�
�Vu�	.�� ������#�2��5ɩ[�����Mڨ���^� ��!-��o��z���k������rI��zH|r�&A�'��;Q�����N���%�~]�j6ͼ�PY�����$�u;9[�XI�&"�~���3k���J1r�V��\y^�
 "�1�'�8��Yf�I����h��߮�q/����fz��������i���6�{f��mU�l%��C:g	��a�R��vFrR ����p��<���of�P�g+_��ȧ�WK��:�K�"-����6�K��ޥ���/U�&��,j�J�L��M2��O��P��4���ڭzA$Uzb��?�� �0�\�[�)mlr���\6%OߊO�v��C�J��#�6�*d�6��-ܢ�D�t#ؕ��;��m���=��|(����[#�ݥ��gP�+�@v�[������3�	�N	���;R��e؎�p`��L��!~��e�Ysߛ�Sn����� �[Y���6}��x���K+�YD�l���mM��~D��7�1`6��Q�z�p)��42��ԟB�b�W bλҾ�F��b�w_�q4�7��y���	����D�'��Zx�n�u�z)t]�ժ��տ�'�c�'9�ĭK*��8g�ىhQ����}�_�L8'�~-׮ϲt�b ���k���Bo-��K�+��|��beu�$��H�Y����F~H�ko�^�%�ފ�g85B���z��R^��?9��#�kQc���u8_d]{�,�^��"|4��i�[�L�=��r��\Z�b;��
z�` ��/Lz�Ϩ��ڱ�]yQh�j�����v����C���	�e�!�˓�v��T6�p�~T�f���N��f��6!�g�?du��;�uS+Q�0�#�f7���gh�C����|u3錷���w����TCж���|�o�l�7�c����k(��ez�>���[&�*G���X�E�"ϗ�}��׻�9�o��9.�T-̣���;Z�K�ǓvA�����}9�#��`T|E�b6do��k��8������#-����C����)R�Ѿ���X�h�i��Q�cψ��9���|O��ͱp�I^<^�C5�}���J�s��>�|��{(�[`��� ���5��pÕ&!x�Z�ӊ��W����!s����ę����o4���0?~�"X� �������^�I��M��a���r���_9h���ۿ��$9͂824�uwȽ�|�$�M�CHB���満 ���.F�����n�+rqm\٬Z�Z0�E<�S�e�-6F͎�y&��ِ���c��QR�U2}�I�`�����y�U�K3l�&�h�yY��8�����Ҫ��o�ϵv��,O�<�)����u7��9M5r���=P��d�Z1��j٤Q���6���e�?ZM����s���8>Q��۰r�~�����j0�3��̀�?�}��R�b�1���sⰒ)Wp�fX-�>�q��b Yޢc���r
�p�6��3f�H$v1�g�E��b���%Y�T���-!$����J�"�`owe�{� ���T��L��u��"#ZGL?,��6z�A2�ǯ��MO��u`<$�c铅PC�J"���#J�m����X�`�xmmXJ�Z����c���&�
�4I���_¼)�)��o6�R9;�E���-��r�$�}2Dt����k�e��^��BO��_o1��9�����g���M$'�x��ɖ���_�)8��K�ȺD��A`���c%�2zD�9�f$�����Zc�lR@b�X �;!�/��؍fo:���q�t�SP�c�a�i��e���ܭ<ϗ��u� x�y�u���K�8�m�����q'-�:��������BGH԰J��c�-��R�/!#��
������kr�ˣ�o�?�*������/@	+����p����-[Ϳ����q~9�Z�`��,�`0U,G�bq��׎��U7�'2w���u�5Z�;��T���-n�Ǹs��Q�)ίH�O��c�*�t��R��ͮ�V�kL�q�*h1�%�-Q}�r�5g�Es�"�_���Q����	�Z*(�U�pF�w�9oo���~�;ޞ���x�ʢ��kWK5�%'��C��G�F!ʜ���O�s1�k�fK�I�:2g>�"i���No�X0�"o���k����(��i}��G��2O�Q���4�2lOn�o�'=bR�T�)>�&��~ ��^8�W7]%nS̙xw�e���*H;�T.�\0QM��/��fsL�>=Ƒ��'�3��҂�<.Q4�3�̚��U�5
��\�:D�击�����x�1�Ū���`���:*Uv��ʗ-�ˌB_JNCAW���Y~�=TZ�Q;WmB ��H$Y�#<���yK���0z_	�~p�Һ�T���ץP<�x	����D3]���^���&>��bSlE����ݏ}��q�{��YL��͡�`����BH;}Z�4=f��^{��zL�S6Kz��6���:���ϊ����/J�o�V�Y���w�.X&��/&r�1��_v	쳨��U5��t��t,��<��6?`��-� ����"����%ON��P2hld-a^C�Nm%�Qb���4.�(�c�2e��
vZ��IJ�[DL��i��#���t��~��Uc4Ѓq�cY�����I�4גe-�W�����x�E�m�M�S���dC�:X��1�
y�&Е�s����2I���ȉ	���0R��F� ڸ�<��u2\N�(��K�5�f���I�z���`�/�Έ��ҏygO��*v ���n���ʅ�T�_~�5��"���Piu���ʶb�ƣy� �]Ҵ�y���pwA�'ī��Q5
=�5�}R�x��/���ajd�gִ��5zeB�J�C�Cl����_h�n����S�Va�X��x�좛�l��R]:�aUz�S¸
���qkX+�`����J�v�W�d��F�4;Z�cޛQld�T_3��+�;ق��m���|WE�	���Ǚ���!%D�
 ���G"�^Eݠ7�N��DM{ϼ7�B-�}��-��´B�:3���$�|���e�%C���HfDz�4�',�n�]���,:���Y������/����q`b������X�S�cA߃��B�
4��7�~�W����ga2� ����^��C��iPA�i�vJL"'"$S�	U�9 ?����G�x��te$U���U�`%/���\��Vݚ�tk��� ��^{�vn�>EyR9����\\���)�\|�kR�J�+[��p�`�D�2{�x���R����)�����u$���!vm��O�}��j���UɄr�$H6��ejA
�Pm9�.y��Ƞ�є�l+`�M"@dЭ����FJ3��A�w��s�Ȣ�:��Ĩw	KW_����R����Vc�}/(�BO�	h�?k�U҈u��`;>w��p