XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_/X���X�Goş��V�֣$�d��%�V^��z��&�=H�D��	&��גۢ��"<�[M8�ga�W<�F]%4v����Y�E����Ђ��čAc9��cﺇ��L�q3p��� �9:@o8!�l���[�Mx`}��U��ů'�t���f�M`��s��d}t=b�^��ҧ�Sh&����Ȍ7/�`��b+���؛x'��i�c=\:��Bzw��ΰ{�;�i]*&h����Sw���U�t�l^��仸�k���FFekwe�"^7�JUX��"�?���+8���S�0���X�Iq��f���!���/�R+YK.�W�p㬗&2���'�&��t��J8rhG}�6�~�d�E�x �(|�h�>�U���b��j�>
�.�<X��T64�����'% ���LJ�l��v�΢i���@�چ�7?ݹ�U��ѭ��Ǩ��@CS���(�r%臬���T�����a�+���-��ܪ�U,���� o�K��h��@�,�=8B?;�8�:��}m�$7W'�1ޡ��Pi^��q�҇Օ񺚃�#���Z��*�ě`����/_�}R:,W��4��f���=w*���`���X��o�ç���*�a�]\��F�=�5}>�
#�֧z�X�Px��,��*��z��E��̰���}uk����5�V��$�" �9��|��B��Xϥ Sz����6��c-P�EJ��<4�$x����Pe�ݍ����	f��fY��鯑7�f���E�X�n$XlxVHYEB    7119    1360�RrӌL�9	W�p		�����&�yCK�Sw�J9=�5^S)g��"\j͈t�'<�����/��IdҰE6��ژ����A��,1�������0���������>cn��XLC(�c|��m0����	�u4�ɊO���Nl�|3�)�NlԽ⻇7�k����V�{���´g��G*�I�ņi{yNY�}�ߚi�fZP��ʣjT@�~�������\9{/�,�!��օ=�Q������]�S�%J�k��8j�UH�5�D��3=.�A���u�p�Z��G��P-�?�dn�$�.1_f's�njp1yc�>�Թ�k�,���8��4>���N3_K6�E݁����Jnf�\�R�$��6
��)�P��R�}�����bN��LWn2Z@�����$@���^�)�9|���2�z;�{գ�*3WS�y���{�,b�W�u��
����l�����Ql{\=zDF��f�\������Q�%��4�k�H!�"�jM�iv(Α $��ތ�#��>���^���֞V�'/7�Ц�q͢���T�δ���L��j��7F7�T^�w���}��$��)P��y�@�r�8���>�	ڸ�y'Y���_��M|��2���aD5S�?5�y|����<���ja�k<���:�m�����Y�Jm�S��������\ܤ�n�BM�3��M݂��|�[�&��{�B�UZ|��4�fn�cr�[��b,�}-�KOW�2���sx���)!�C/&E�*_����t�ߢb��Ψ��?�1͟`[����;�yc�޳ɝ��I�`�c�
���9�:�=�5"�ԓʞI~�Uf|!e�*�0�恪|lGT�@s�]![����} 7q��R	U����� UVt7�kW��#�b�� �� [#��*11��3!�bA�xz��u�����0_9��<��;֯T�_�6
&�����G��܊��H�8�6��Xዣ��+A��3���
����zb�-0�ɇn�c���h]�i�dqE�_v�E@y�0861L{pdY�֎�(W2~��^�YF�j�0߾�>{6�%*��M����L��\�ACś���F5��B���FiZ��6�9_�H�U���D_�ɵ%*&~�/�.���8z�6����r��b��S��ʡ�/�d��\3��z�;��`c�1Vr4��qa]�^��A���~�&�6�p��DRp����P��?�l�o�" ���5o����]ZB�|i��&��用����~�!�1^(1��(���>M_����hy�GPUf	�H��ݸ�B]ͅBy�}*�*�xO�Pݻ��.2_��XB)���)d^<�KoD�7-fߖ�T��@�_�;[7Q��)F�h�!f9"���	oA��O�g�i�Siβ1�I�?z޹�e�Q���j#����]il��U���q*�tN&�έ�A(T	����Qm%�^��2�L-|m�/�{�<&����[�9�Q>��~�p�˥���ve�Hfzp�H_UH+
�ٴD�6^%�d�GUc�����eBrD�TQ5>|�І�0�O�kօ~FNX����D8��N*�=��-8m 
��g�8�Ï��Q��=P]�rW}�
QL�3�����S,:���D����v��:1�����@;�����J�8����X�[�`�[R�LTE�\>��p�F8ݳ�`�L �Sߢ�W0��2$�I��.��}y�O+(�1Όw�O/��s}�d}@T�&!k��҉��Si����2cμG��̿�"���\����vS�pڡ����S�v�ys7�,��K�mXT��p�tz�b���
��`ry�1/?R�g[�a��8b���	�S3�KN����df��Q��b�l+���� 
t|��fxŵ�ϰ�j��Ժ�}����Y"$^��
��\?R��	u�S:{,���S<�rM3<���������'j����^�^�G�ެ�����쁡�B�������]��i����C�f�XwI����L�!.�ش�r9��|�?Qo�sA�X��M�69ow��2p&kBO�͆�����n
��E?&R;廌̆CnjS�݀�D.D����48Gq�%���^���7>4�S�W\�;;�9�ք����q��G(Z	t��Ddw�/��7'�k=�1�*s	O��YCE2F��ο�W"WP��A�`6�R�.��L�7rpg@Ԩ��6��Bm��x]h�.׸�U�:*���I�U	'/`3*��� � r=J��9"�)�o^o����EM���yqL�����tK2(���,$��f�me�݊���B���Fu�|絘=��9�֘b�?��hco�?C��a��&)5��z���D1�"�U\�CFmn���?S��S��c(�d%Q|O�a�)�c
�pKh���c����b���Ù�����9�2�0�����v~�[lC-ᔡ�>�'C��Hn*K�룣ͤK�� D��	���mb̴Mݲ@On���NM7d?�h8��?�dГ��y�����X��2�����ޥ�F9��k2K���p9����U����T��ui܃7�]��gU>�79������u'Q^�!i�M�;s|`z�������}~X%�zkʗ7��F{�[��ヅ�\��:Ű%��%����p�藁�nʝ@\�y��euwp�e��'�$ǁ��=��,�V�E����X��Mm<Uᮕ����;�^�'��a��3��ȸ̳C��cs+,���|݉
��,%�|�'�`v9�L
,���N���BT�s*|�G�<1��Ug)ݓ��~���4KC�5���c�aZG1��]U~���z��=c�¯�d}�u�AJl�]�)	��j|��{#�5P�I��O��:�����/��֣��ʑ������>�=�}��i5����òb檸���!5��c���s���_�M8�ȤZ�oYG�i׸�0���j�P�Ț��-���i�L�Ut�-��/�0=��~��'����L�VA����E��Eb�tRb@�rkɦ��p���ʞx���	C���u�_Q��/�/��@���]>�H�G��Le��E�����~����K桇cl��٤�D�βZ���Y��>��(X�:oUȟ\�ޗYk��1��t��J,/(0*���Kb��V�O�Dmy	[$ ��B��d#'�J�y�~Fwq�@O���-�ϕ�eazt��70�P�P��J�� &ut�6�7NT��؟��1�v;���Ԗa���dЮ�C�D@}jWP6�8eX�1�᫿Jp(ا��A��z�/"���-J�b�$�t�A�m�rD1���&m;��w#�D
	�}���r�Z|��Xs`���Zٝ�Ǡ#_˵#7	%���pv5/8F�G�ח]"��0.��A��+ʨ�em�����(��}�8g�3��w�V�'�7�I�-IQ5�^�8!fx����i�5���<��<�zS���g���|�8��ä����ozQ5^H�L�Q/JG��Ap�'���#�"�R*�)���O����6��/�i��R�!E88����<?�B����x�j�v=!�mLА��s�1�j��fKN�����
�_7l4����o=��gP�x!EgHw�˶t� y�+��%=�x�5�� �A,J��?>3���>eUQ�r�[���:Ɗ�!��x¯��0X]�?hU�Œ1��_���O��f�����1��d��T�9��rCDH�S�@�@���2I���`�#�k�d��@X�L#-:5O:(/��,q���r1�̎o�*߻�@����C��W��(�{�g�`��D��	��>��%��A��w�i]��[Ǔ�)ۏ����9��7y�*��<7�D:頺�� yvt`%�EI��Dˑ{殪�T���Q��2I�wN�y7���⭞��3��A*V~O<m�(�c�׷�6��1�1�3��H�s��K�r�{��!RW�����e��v��K��A*��ȑ����i� ��[-����Ӎ�X���	}3���.0W�5��p]��YRiK�Fd��2~�[�	�ݍ�u�7�(���ο�t�&P� �8=�?$��)?�rk��C�2��KH ��фl���F������,԰"�?.�0 W/~���:,(���짇Ӕ�uy�|��k�<W����cF�z*݂�u�rfѯ��R��?r�;k�7Hϣ·�4����#��<���|�&��bޘd���$�`��'n�v���A6�2~��eO�l	M5�B6���F��{��8M�̙|���۟��Fl���@��r��X���p�я|e�����_Wv$m~!�=w�*�����"�⣴��ʺ����Ɏ�Gҍ���E��I"I�u,u�&&CaYhMg����"�l�����f�*�|&j&{�&.��r�m�-�t�+WS-�Z�(��K�V�>�������
|�b���NfN�M�w�sٯ)BkQ��� u���D']���	��.��݀�
w�����L�%Nm��Vq���\~j�8Y���Zz!(�ar�z��c-�K���yP..���y�&s.�n7x�D��!�ҲrN����X��>̚�ӉX�3�����W���f_L8��%����������E�Ű��A���m��~��SO8�����^�;{a��B�ɓ�k�O���QN�ž`�]��G`3.�	$5TD1Pj/AgO�C�g �j�����5���U������9�R%2o�=����S)�0I�Vicać�Nma9G��ZL�k{mY�4��7���˞�l��/*ϑ����`*���y�f��IKC+βc��%�7�Mg�����J���~���9�g[b/O�'���*4�|'r �P��0��J�&�Sd[��FH:G$�R��ƻ����s����x