XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<-����X�s���ϒ�If������\M����
̈́Η����o�e�Ȓ�4�%G�ޑ�k#�M�N�<�����~U�Z��?y����S���3��K�����\�k��ڋ�,�ț���R�*j��=��4C��3B=wO��.�:��ǀ�B��s�_
S�)R]s����o��\������<T�aV���+��!�?~.�zl+ϕ�v���y ���-���H�#�and`����6���Ԭ�[$���7��RS����13����Y
3��)�,C�w��8��49N��m�]��4'�Q����h�H��9�f5�?�����?�\����œ��;��z�d-�3��������ҰC���:d�%%�+3<�W�䁨�a2�x��/�����MhL�(�΅�Q��0k�{TЬ�~�k��L`'? �ؠH�����
��U�<T���x��j{m0�$�X���������u$��C��ф�Ǖ�x�/T�zt�N�CP�~����W��5ڇ���z�)^�4�;GK1�Z�Ȑ?��́d �t�G��K�ރ|u�^�I���� �j�ϴsCE�)M��!��B�X̩�[Ѯx����3N#����.���%厃tP���]�V�Ǌx�?�����kя��,�_��G�R�$�3��Bp3�;���2�{��� ��>#?���L>�{Zxa˖�Kt�Q�["0�l"��-�l�>���P0y�(�BCE��b�����E���h;F�N<9�oXlxVHYEB    3daa     a80�2�Z?���b`_���{ȵnm�6�G�O��.�B��uY���T�{�@�{2,�!il�D[+����̙4A�9G���i����Ģ���o�Z���ヽ*�a�@�Y��H�sy�٬��6���,��V�TqLU�&>_5t�Q7S۫�0�Su��M��L�O7t�3n\Gz��~B�P�4��@���o�H|�e�|s�)F�J^�	1�3��;(++�W�BM�شҌC�E���4g�T4�����9�W��-��I$5Ip�H�W�y�ٳ"��N���}"~wGtT(��(e��3Xq�屬��ᚚ?��W�:׊�$a��4�԰�$_��G��7^���KU���h�K*
���`5���5B��g�v��zb9��������\
:��A���?Q8l� ���@xw�����0�{=�Xʏ O>�R��잏*������7�']y#߃q@�`���(j�ԁ�żʾ>B[9�����L��n�>�M�h���Ƒ���sS1k��y{�� �y�>d�i���p�z��z΁�cM'��m��+)���P������]v��R��j�T0M�csʡ�<Z&��K��f�d;f����V�A8�S��q1�F}����_R�H��\C���$�Ԑ���uP)���wO뀡h�Zp��]�xpd{�4W/:Lp���s�Z��n�_f	�D������}���y�#�uo�d�GW�M��x$A=B����	 @b�t�% j|�~��TH�kM�)�z�<�5��u2�w?tp��*~a5��kK�|��{�W:���D�3Wk!g�߂�؃����2�Qd�/�y+�\���!���n�[7%5�J����ڲ�FGv�>�\�=員mG�~����D�,;R;�cx��P��=!T���;Ww��+�drP�����6�9 ���$*��?��U�a��+�W%�p0���u����i:z�:���?fn�T�Bh�]����^ڎ}���Z�t>�x�l���r�ZQKK[ ��˗: x��R��"���'[��@I�e����������T]��7FZ��|�|C&i9��"��ѧ�wA�~��q������|xϫ��yr{�s�X����/={�ʀN1��4�];*��R�����i��":^9��5�?QĪ���2xah�"r6p�]�i��f~Y��O�S� �'\�vR��%}P _� ��]�]Y.2��hl���xb���	��3c�tH��VBN��:끯�w :���V$�XZ�nx8)&c Sj�LZ�����IV��۳Z��}x:qć	R�����|�r��w���M%�S�b��lǫ�mŬ�X�ܷ��q���z&�������/��d�����)�����d~�F�eޔQ��YF����_zG�� �E#�t�б<����	��o�������&0��,7�Q#U�/3�ի��{���r4��(�[v�E��7�%U�a�z�J	!^���yQ8�F�%�8+R����T��x���(1?q`����~���]��������sӭZ��Z��D���7����;�\-8�UML<io�3��w���l���j�6����}���@j�f�D������w�6��@W�FϪ���Bb�@|� [���l0y��F���=dS��nU�W�eC���b�h�LG5��c�ƺ����`���|L/I�)岓���o�G�ZWȪ�(�ke	۾o�H��ե�܇�1;���Ч�����00�#��c�*�(dϻ�ʬ�T���X�d|�S���[��H!4���7I�x�5����_�I���R J�`Z�>~M�>Q�s45�bs�o��`�쐷����ʿJ�d!�%(�g���׀|��?d�����E��U��b����\7�T���[���A�r�ӺT4��NQ�w�����#��T�J�!�?K'I��n�������F@�bFn�w��I/�AE��.���{}�A�%|V�%�p�} v%G|�?���;��妠�ӣ��5P� �[D�8��
|���螏D~/¤��1�u�ɲ�0�ؖL���IE;, �g�¤@��;�K�V������ ��/��]J0@�;*w��M���ZܤTa@�?.�����:&Ns�����,�  �=M�B8N5�\<�����jTJ��,��{�� �W9�%�B
\�bH9���J<�"viP�Ô�q�爕k�$�'&CM
�C�-<dsc��T�*�P�M����iԬ ���GD�	;+�r�[�<O0�L�-1��+'m��?�����ngc�r�!�5$��k�q]@;���;<�'+=_4O�QF�#�mH����ʅ����$�g;�٤��g�C�փ�nr�zK��T����1�FdT�O�kP$k<lk1�|��c� fT�6ci��'c&Q�����(�&q/͐_��.zE���Ј�XL���m<��o��j��R�1~Q���6�d�.45"��3�V�k�Sl<�D�����xt���LL��uN+	�ʡ�ädb�H�|4ĺ���m|�U�ϣ��	�����U��h?�i��V�K��#�V�̧��d�V��ޝU91�"��w��Ν���J.IxƷ���z	�uX4��ϕ?艢��x���,��;�Wz>�_Y�