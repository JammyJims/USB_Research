XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�	s��C	���#���w3N�9!�IY�'�>]~1����z��j�~o�7�J�<(!�g�)����.����¹�/��q��fQ`O�e����.Z�%U&������o�^ʷ�2Xm-�|����%���&������Jɉ�Ӈp�V�&��G&(�A���z(B_B�֙�����im�pD��܏uU�n�{@SU b��8�"s���*\�{�;L�(ω>�F�=��m	m-?:n�`vn�U�-I{��J�z���E��ϥ��=7�~�te_f�RZ��
'9�p��J�'}���EC8�`��Y�j-������(�>g�;�w �nד *�NW���lz"�+is��5�e*�e��=��O`,��Č����ƨO�W���e#��mw�Q��.J�>���z%�C<rE��e��9��:�w���qq�ۀw��n.�k*�*�)47��dq�]D�kk��F�����������j��_��r>�����IDץ.Rl��[.?&��r��(@���,J�z���+&M����
Z�Cd?�D�ZtS�3~�ԗ�T�`X�p����P:IR�\a��Q���w���卍���F����]��Q�m��d�4$�~��B��&R5��ʍB��=r�.�~}
Ҳ����l�mϷ`]d�L���B�;i8tP��'M���M�5�a�T}w��;$+R�j�|�C\�[��sȈ;���e��s"���q��cfp�w8)1嶻2����XlxVHYEB    2d65     b60����e�yFx}�Y����ƶ��2ߜ�vs��e�:Ʋ�M�D��ٍ���T�U��V���k�ldې7��t�s�zo4�`t �{j��w��P��v��/s��T��I����I6'�ױD����aB?L�)���$$�V�<:X8��*���D�XVx�h|	��a]��S�rv��ԃ���#��!��8i�g-�?!&�)���1�(kXס3r�y|`��d�ׇ�g;~�+�� ����tB��(p��@���qk�롻�P�s�<ǹ"��E�v�$�) �+���1�f��[QHJLr0ڴ�i/9�/0���9(Wם�qG�ZO��nv鶅Z�M[�1y��@��D��5��Ʀ�>�/�_�}w'c&�"G�+Q<����Sc���g镀���P<Q�4(�R��J�e� ��VC�v�ȉ1�~�����N�.��t2��KyV�锶W�$�#�.��´'����;�k� =uf�}��RI�8WItO�P�#~��b\�=�60<+�N�Ă�'�ʭ�r�.�0}��� }��eW�op2���_� @�9�5RMj��Ͻ��G읏��|�&����t�i�O{"�G���m�;�i�kU:t�������4H>'*e���3�� ��@y#�����	��xs����B׍�p�K�'���q�ߦ��7a��B��\A]p��3 "p�9��KmsAd}z�c҉�e-G��ބ���c�W:Hz���!c *���K�!Hi�	�k0�=����C Y�0oWt��ƞ�Cℴ��D|��S����w������ǧ"g_������q�L� y ��$�0P����Wóbn��e�A�@|5�a]򘦹'@[�$ſh����?��͢�����m�ڨ���UȩE2�!�B
湫t�oT��g�.z��\h��Y���C���K�wh ����YO�R�6߅�2^���2��3<0=�w�:�ڿ�4��`�ņR���
d���s$I��w�klT<Hd��A�К�����dI	��q���k�����%���urg�RαY�޳N��,��qS�� �Xh �Ƹn���_L֬0.P��q/*����E��+M%E�YGj�~�b�{{f#@�[�[ӊNp罁��"�!�&����d��6Ǻ)���㈛D&[����T�W?$WOԺE�Q�Q6T�������2�:�Hټ6�'RvgA�{���y%��%�T�R?�s�|6[�	��4���(����� �m����r�챱�l�(˰U��xAԕ�FF��kx"��i�w0����<�R�<�x��E��q�ֽ3�g�����ѫH�Z?Oh��E%��D���u���������C��Z�1;��W�)T�q,_t�(�u���п��E^�+�.�Ñ ���|�.��-����գ�~^I�ę;��D��aV�;x��󪁼���W�$��f�xh��(�t�W��X����+M��+�]st����ý߇?Vq�����^j��<������J�'\�q�;b�z�]�w�_l��k����*J�X���~z���Ε;�D��G��j���E�_��l�O�A	�O��LD@�Tv3�1�چF�d�'f����˓v�"�W{���toӱ���+�( M����KD��C2~�p��S��
/�V�O��2���3��c���ᇍM�S��̝^�=�|ٴS۝�.��6X��f���Es����o!$h}�Q������.?Re8���	/��N�e/wws�r8��\Li�q��a�޴���)�cOEz_�ޔ��6�s��G���ōT0a��AZ.�~�G�",���=C'��z/�muV렚gڔ�6@zb��,������fq�-��u��Q^��M``BE�Q𧻚�-�8������po&���+>������n�_�.��u���_�V�;J�	�!�YՙL��+����Y�CQ	��-�"����,�\L'��AM�`��4&A=�����E<�\�Zٌ_}�C����p1<�v� ���,U���ȑ�j쫀1y���&v�\� -�r�X�5g��(�F"&9���C�Z��riϙ����>�[0�|��,s�g�f�w�G^�D�f�Kt�E��c*6$d� {}+^%6�_�6�y��iZ��?��R�S8{͢U�K��=� RD�j(�2R\�C6M|fՠ�C�5�~N���I�������3�HN�������������N�ү���aw�Vʷ�j8��k33�~�lm���^F-u���T��h�SY��N�b�)�����,�<gnX�I?;A�O١r��1�D&&���k��G>���Q:�w�?�|��J���"�P	��I��]�ؖ�	�����bXQ&Y6���Hp�[P�#�B����*[*������4(�pP���y�M����ƕ70��&�m�I�#]Y/fцp��2��Đe�_�H;�*;�`�W!��t�Kz�O;}���wi�>��[�*�գ�:;[�f�W$��k㹄su�l�]ie���u�:�L@�P���́���WU��7,�� �~o���MI̓{� <��4�m�^���a?��������HdIFE�XxP�|[��Y�B\9�"�1�_�\af��G���1��/�`� �t ����;�G����L/#�t�,YRb[?�lNۢ�s[��"���#b�y�:^�՛�i"]�j�Ӕ4��q&��In]D�RkL�?4��M�AD�q5{�'�1&|)r�ҧ**��4PN#��;-�-��&�dp�"
�p#~+�Ҋ�7��Fm�[��G�g8�ߢF��d�sj�Q�(RXL���