XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���K�
l��t�$b�]>)��'���r!��7�WT
q�@� )�9��ދ�JD��"iU;j�&*oN���t[3T>���ֿK���qBI�jrEE99b�V�2J#p1#X�"Uv�R4c��fz	��)�L	�9ؐ^qr���nj��n<\(h,&�J2 ��f8j��� ~#؁��
P�C!8pAA���;c&f�c�jD�?V>�H߂�����{lz0�v��K z~	��Re��t��[ԗ�m��a�,�Ȗ����#�yKR��ZBD�����������W��_��FU�8�Ć��1�%@�MZ7�H���l�%u�vC���`�d���"^�}���MĢa��Ҷ�>�
4��䝹�V;�UwVY�h��'�����3k]s������~x��6i���?�S�V�v �"�%'"g��}���#oD't�*R����
0F�M��y��(�)�
���pc�*��I�U�
Z�*��՘6t7Wu�<���Rl�R�6=	�hA&�<�2�rE�VL?��[����Mϑ!̯D��XQ3D�?9��is)�+p}����)XA��>UJhw��<Z�������5�{]�ɝ�5�*Z(�#�OIr���.}� "��#�,L����.����p	�e����8 >yWMK��e��&)I/۽�����=���Mb��|n�A}�%)���C�Sd������f����g�J�c�X��UX	9f@0=m�ņ�5��.饍�u �cXlxVHYEB    252b     d00�u]x6jRxY����y(r�A������w ������EDS�1�-հ����,��7���U��{����-��/R�wk���͢���Y��X���N��#bY�ˍ%�w���"R���Ww��t�ٵLW�MRJQ���+�0 ��d��V�o�mI�~3q�:{�	P|8?^R�Ƴ
S`����ki��=Uw&`��	Uss!��ZIA �la)�0��E�A�o)����S|i�k���9��q<s_>TF��ʬ$��7x�������J�o!��>�������>��_�Ȟqu�C���?J��B�����;��im��
P�$�A�j�)ėE���}��E��K'�>��_�=��!w��&�B!��+�?�2b
O�1!�Ը\T�����Fsj6�K6����1Bcڈs��{+���/L��#�μ��X�d��m��!���yIڡ��leL��?$i���G�yU�\ȩ�8�Dp�|d<�������a6�)�-k��T[n���PKX�nB2�]�0��Vl�(Cl�H�v)Y�����2P�=���NX�w�g���ه�铢�|��s�~�i\�c�%��=�ں�;aD�:���qv��EX����yۉ��
&���Ru`F��Y��zE�(=q4f�砙�f:��l���S�����v̜~��z�2>
���|�躆�U�m�^k˖L�>}Qn�EFA�V��CIug�]�a�=�1!+�W�h��!��3jܥ��K0����7�VV<�;ӊ�{hN�|�W�]���cՃ!�Š'��w��������ݪ7��`�5��{��&3@+Z-ao.᝵C-pYaJ�vikJ���\�I0'�#�í���N�S�Lb�9��w�3EO����Cqq�~��G����Tno���$>`� �����9.����3p�iGHv4���Q�u�I�v���u��4h2ɴ5ji��$k_�x{�ŋ�^��by��,�m]{66˷�߮�Gփޑ�����^QB@|�0��2Z^ؙe����y�@�yd�Z7B�ByGq*,��OB�W���"(���%�����!�n���kNҫ}�'�����~����v��^�|�S��ߺ��L��4��,@I�B�h�
ik\BZ��=n�yp�**O����݄Q��/�fp���~Ȅhw��v녉i�V ���ǭf5�S�8z�
J�c���-ز�����Q�%ќ�� [��M�����>k1i�}^�	/3"�eF������ͮQ��N�����8+� \ٻF����o	���B�L�Ӕ�q��l���PC���-��<��~#=HV�r,��ª�^����V">�>ira�N�᨝�.�rE�Xܛ����x����S*��݈�2đImw3k���Z�?ڬ�*53�U;��?�X����\�����[��l_�wq[���Ĩ洠�,݁�~��h[ ��8��DN��
P*�ş�V_�1�����mQ�D��T���c���Zj���Cе������7�b�1;d<?���*�t1�H� '7F��@��f�t� ��>�j���g;v�g�V� �y���%�6w�t�;/F@T�Ս�sd���ť��R��}�'ٶj>.Ϙj�"�jΕ���tj�6Z>��WNrQgU��j@��9�ߠ��f�m
Rj���+�l��\:�2�$sU� Wj�D;縀��>���2���|�믞)�'��.�K�s1���HP͂S3פ�ñf�1í�XL(8�t��:�v��Z���`�x��"�j�|�c�wvlQ|O'9{�������j���Z��?Z  1__%6��?M����D�d�;�[�k.���ו_���2ULR3V���V �[��c��h�e�8��\�*�+�]лwq������_���u�x�f�	W�NǮ�y�+p��_�����P��;�ؾ�԰.�f�n�]m�/����V���I�����WX�X�5���A��v�li�S)����6"�&�G'.�)9ZUXZ0�_$L�!P}��98�<�҆_�οbwEy:��p��B��Ep|��D��MxU�	�g��&�-0b�|��*;�J�7b(�g��խb��]U���r"��C������+�-�2vq(�M�M�)����fԏ3�>�1!��fw��	4=��!���W�KȰf��t2�ws��kg��!�J��VY��a�V�KS�e�g�K4/�S32�3�����נ���C���QDy3CB�,��~F�,K�O�x��Sj����;Xg�ÿ�5�K\8�>��J,c��#e��nR�I��P�f`�l�ڕ�D&�q���u2����5�v9�r�� ��E[!������^ve�r��*��<���%�L7X�4atY��-Ȥ̍��=�z�oF��ې�[	W�#�z�>J�����)ņ�e@���	���6���J;��V�=�_v"sI�[� ���G ec��ɏ���� Ĥ���3�W>}�7jY��\U���m�ܩ��t$���|}�@ �3��w���MI��X�cD�"�����x�=�A,8�V5�Y�ݶL,<<�rO�1��o�
���ܯq${�{��2��P{7��+�I�x��RvS��b�_M�5a����f�󊷔�>���`�$���W�����޺7°@l`|��,%H������T�����\��;�eUҺ���_��Q+n]>8����b�h�\��z�q�\^�R �u�,řw i$cyh`ćr���Sۀ`�|�7®�_��9��ݙ��~Qzo�e�\�4�e�X�#��E�ϱ��X��:�tJ����3��.�	���Ur������Z�75�[[�3$����Ū"��F��籥�Y=�G�M�G�փ��@-;"6h�aڌ�y����Y��0;��9p�Z��k�^ߎ�*B�9Y=\���3����/��Q3�Ĺ�(��w��q�5���ۀ��oqH���6���� Z�d�Pkp�
ϒ�V-7��	ɸ,���Zj�~�I�����q7�v��㎿����;��q;Eߣ@k ��>���+� m�o7,{��٦��կ�z�Ғ�Mʧ�$΄�u�n�7���/�i��ƺ�8��D <��*�|Q�g�E�:݄M�OA��!�ukPN�-dn��g�R)xl�
�)N�iğ�g�{�}�\��qK%��v�kGGy��_��$BҎ���d+�~#�ԵZWO�Â�t��4���^�h��B���2��0G�.�G־>��2g�+s�WM�x���X��G�+7r�|ޣ�qs������