XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ʋ���zy��x@�����wq,���R�(��]�.{V{ ܜ����E�<k��Q@�ir�V�X��h�^*���UQ�ȡ�;�Nv�/�7�P��]{ӫM}�hk��
��ӡ�å_�b"��d�d��"q�4ܳ��`�?��(��G�?ExA�28���r�(;�߲JƊ�!P�{�8	I��zL��	�1M�F�,%5�3�b�T�>�]F2l�e�aU'��p�v<�lL�
e$9���g��[�T+�P�	�W�G�U��p^ы$�g����,�X�.�-�-� �{%J=E�2�ʊ��Rʧ5���ß�3���C|��R/��ƚ4@|���w�Yu�|X�BN$��j@�|Ha�&��x��Hwz��r���1�@���C��j}��Fk�6���^�>�`hB� a�6�	.[\Tw���������Gt��W������?�{r���t.m�TW_��^�y�
���Sж-�v}�@+e�FZ�*�:OD}�"���gn2R��nV��>ӣ��?,�?�(����.���Q�{
�Q��^V�,:=h�I��r^�cc���xd@t��y6����V2<J�I5���Z�����.KQJ����/Z�b�y����-��.���L�LEe���0�-FW
�ړ]�K 4�TZ�m�����h���_�@�/8�9V�Ԉ>�3y[NT,��vU�{�H	����k@d�ȳN8��z�<�U�g�zz��,�[�Q9}�k��)}�XlxVHYEB    1849     9f0��ׅ��_s�O�^Ѝs�\f�eJr%*�
`��Yf�ؕ3&�g�������S~7vK�&S�#,Y���B��pJ��&��o�Ch�G@����ySl��D������xи=�-T�����p�Nű=	F"ށ�� ��J���=��Y>OU8'ɺA���󔚦�0��4��T���vċt��A$����ة�.o��F�ѭ����C&�f�:/[ǣ��7��^�s:����d���Ըql�a��Q��%[&Q
����S���������!�i�"�⶧a��;�ơ_�����,ŉ�D����l��J:aXc0���I[W�c�Y3j�~[b�c�fO���tSC��M�̬z
$n�Fg���Y�ܮ�**|��l	c���7�<p֧�;{c���t��S�L���w�E�t6�t�(h�z7)��&�tg��k0�.��$t���)0��_fg.���/��H;���QKؗ���fO�@Jn�(��0��W�67�P�o�$�Π�W',��<,oN{����y�z+v���C�����#!�J���e��N�����O��{ �\��_�D?��4�(��-/�l�Ю�ɁV�.����<��a���+��W�7����^�����ʖ����wc�eZ�O��hKT�\dq�x"�2WN\��9��x�T�F��l�d/ �� �?��&�=�d+G�N웸�F��١�u�d�ӎ�#\sVY~�Fl�[M,�%�y�)ȓ����FvSD�mB���e�/sy��xo�v��6	MK&L9��I��>K�x��'W"�o�f�9�0� �^>l��p�|��*��i�G���}_SLt g����ZE/h��xe]��kZ��rǷ�1���g�L�ط��c)Kxz���܄�����i��k2eT^A� TSm
�3�Sݟ���0(�����)�ֵ�Fv��w��$"���ܗā�žD��Ȏ�X���<�R����c��׿뫃?�3x:~\_��G;zN��Ɨ�tV�q�'�l�N���3EfӖ�8�:#����nܵ�ng��ql�����4-�y���Kw����2��X��UՐ}�ȱ@#LT���d��~ %<�h�#�w�`\j^/1|�4Tv����˙VYGX��M����nZ�tC.\���o��t��B/�s˅��)�u����m�= f�$ ��S�BW𸩭��D}*�m��+w���Z{�Ty�sn�[��!x���-�f��$c��P�9}�!e�mqm�oT�v��K�ъ�>l�j�Z�H̼�ڤu>���[�Q0S���r��Z��w�Z�\/�R;�� ��������F��/�5W;��$�x[����=H�	�0tEм��	�k�'m�;�e�/`�p��~Rj�kk��u����_5�)U?90|�����(
,o�n��q�8���)D9�2�����O�,4t���5]�)�p͉�A��Qt�̹�{,3ZE}�*�X�/h?2��4� ��p2e~
��Wž̽�E�(�V4&�4grP�hI��MM���ܬ͔
��3�%��e���}�8,�-���u��[�-g�8OV�u�k{��bV����H��8KD�Fj|���r��2���H�K�@
	����3p]�-�rWmuЩZ�����?L�Ň�t!� !eUw�:#�J6g��Kԫ�g�����)�g~�e-+a�.O$�0o^a߅��zБ,�v?ԟ��~�ϐ��N�Ͻ<rlK�\X���=���R���Q�Y]d��b)�'Ly��EO�o�M̍��KjM�I@n��}��d]�ů���^�dP��}�s W8s	`|����SC��=�txR� a��H�n������ʙ���u�{����>��	���)�~ym���J��2I�[��"�5��t����TB���ؚ���a8:v�!4 PhyȪ6nX���;O�BsJ����E�����.!����[vqR�QI��<o��	{K;>Q?�J�s4S������y�_����&�RJD>֟��W��Vo��� QF
�E�g-%@v5A��Kf�V���&�D����\�� F)R ����LA�\D�����$9�MC[a�����l�t"v�v����3�PX0�͏��Q^����\ڒ�ń�L��B����O��<3 }��:��˨&2�w�ѠNN�� Hm=yg1�g�7d�nc ;`t��eQ�d��)�R7�#�e`��yϢV����g����T/��99L�XiX'���9�8:q�Y�y�
���x@�������N��0�O�/�Kh�V����.��T�S k��g�xP����C	ŻjF2�]���7�`ʪ�Ѝ��n�	\%Q�sƥ��r^��H���>_G|k�]m�D;٦f�xѽ�+�}Wb�*��ƍ�� �G���1��V[�g���ϑϐ�r����A��"��߾;���.�["g82=�y�j��b���N��)X%8Ď��pg�;��'�&ۖ�Y��wFM���K