XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!m��l0&Ҩ�9��� ��_S�#��-��)R��Y=��6��:փbGO;˓xui���A5�mM/�93v^B���O��l��Y��__,�c���k�c�У���[�@[{� +T^'���QR��ʩʡ(�����`��W�������,�N��<�>,��'㲕*�[Z5���`�C����\�~T�<�6��d�L�{��w��+|����m�q�<KC~����ڈ��I��2t��)O��X��,�7:�{��E���D ���
 ����Ho�XS�d,���dO����,����}:Z�W����p��T����c=?���J�`F7h�*W�3c���m�_V����^��/�@"�e�����?�9<ͪ����{������R���^w�/������)G��.�ZĬz�.�Q�m�� �U����8�#�Q���]H����j�ǎ)��r��V�'�΁]�-�q�="�ħ_jW�
_�����5��Q8�f��!��/怞�i0!	�Q��k�+La��<� ����^;�8��t8A���f?���j�A����x����ZΘ���lh�լJ���q&��Q�b�H�[��h#�WckZ�#��m���Q�
`�W�ӝ'��}�,hjp4O1G�
́�v���L�?�9V�Y�R?��DL*��rB��R�06��+�8Q��>��Qm/޸�����4�U�;��s���<�=��3&#gj0�7�žyS�'���ܐ�W�ٜ�H\sʣ�����k?���XlxVHYEB    fa00    2db0����b�T����#�Cӭ�f8כ2��RL���>��K���%M��7���|�����.2�8����FH�Lѷ�Y T 
J��IF��Oݘ�VIߩ��X!VY-���l>X,�(A9�2K6����=��^�s�q��J����j�9�YW���CsM�x���N>k�=�5tϔ��@#җ�INҋ�6�ǡ�M{ixf��^ Zce$��x�{Y�Rv�	c�t�Pm��z�4�z=�e���⬡Fh�����1{Q�7y�5K��swB��c��npF5��We��I*p�U�c�P�*�\��TB�;uu�Z;k`f-�J��#�D,9fi�i{Rc�ă�mL�2�۔�0��B����9W��c���3��قEy��;����V�ϣ�����_1!Y�q��'jC���Ǳ{���8����F��ȱWt%lԒL���薨<a0����v&:*���7�Ԭ�y���u��|� M. F+��8)��9�zٗ����rpn$�`ԊF�����G�H*J!܇;A�c@��ŗ���m���������ro#����1�m{E
�9��#��x�)�T���q���e�7r�BK$K��D����x�ҏ��ᴪ��я�:_�"�P�md�6�����[���+C�u4$�cs�!�O��<_�*r�'ZTn��B�1�!�2��P�69
��L���N�(���J(�_��D�g��%A��%�{.���1r��i�ܧD�w�����[�z_y��ր�*��c��d�QGǳ� ^ �;mX�R����VJ����C`<~��o�6J��9�dn�<O�Pf�7�+*N�!�~L_�%^P��J��0���3��ϭ�č�N��t�;���3ܝ�Dx��Iw�[.oX�#�v4�Dq49�x�v�m�Pa�!������Ĭ�j/��o��}^��3��4��B
�3{nP� ��T���[��	��{Z=�:��Vs�g�i�2"������E�52R��GG�����[�dR��K9:�}�%��9�UӀ�*2�Wp0�)���miDN����
*c�՗���>vy&�	5�0QNe�i�q�+��Z79��;�����M@Oa�}8A��呺��$<
mQ<V`���es��S]���E����Kk�e�f���HԹ�$J)�Y����
��Df�U>[�S�N�������qʸ٭�.'ygk1�K�k�ev<F,�tS�-~�Z���m��$��˕kʵڶ��|�TŰ�V>o���u��M(<��@5U�;s�_T͢*x+���~�������I�Ft��/���.hl��xlb����k(�S��䭾�<���1r�w�������.6F�Y^���v�����gϨW���@S�ަ��ۏY��I��:�� ^����aW ���$�Ե$�=����pI��G@E{�p��j�B��uY��+D,��C���-��_�;	�%J���P��w��p+��g'#DU������{��!`�C|q�ݫe8���j�1�1�bk�Y��k_�3Sn6��Lhff�Mk ��Kؑ�GF�!YQљ�ZcI�cS�]��������kL�K�}�¿�8��������}��6��Ry���d��b@j�!&���űÆI�i`o���"5�FL���!��PZ�tx�a#��c+kVd�Ύ4�����hs��S_ �X������{cp��j%��*�4�Ts�Z(t����ocI���`��]�:P<˪��o��S��FY<F.���o�8��� ��:1}�J���I2n`뷫>Oĥ�ݝ+m��Z�k!rf�櫤1��K�X��V�h;k]>��<�G�<8ȁue^	��]����/�ax�=��F������P���83�6E+�;����8�ey{��Ԋ8YgQ��&_H�G��*6��E���Yo��V�?�'[Sׅ�n���%��8�a�@��Ft�}F�򮮃�+�H��/yS�w���UU�/�$A��T`�zV�3Jhn�Л#H�ܴ����:�.j����=���:���x�`�B4��
j"&''���c�&-��C�)(�4�m,�h���~�"�л�X�$@zA֖T��y��t��`������cˏـ=Sm��-�ES��6�8�>J����;@H���b0xcD�}��7��f���NVX`rS�s�4��RH�pn�s\�H�1�B�]纛���J�V�wT�[Q�G���c����qʘ��C�0������/��Wb��>r�E�l(�ik��­��vs�g�O�_Ü�:?��ʙ�<�*l��b���2M�֫9d�K[�o�px����\W:����̯��f$�?�8WP܈�B;}5X�9��j�T�i���g3�����+����%�	
�������2}����ß�h�W��:���>�����-���P #$�J	d��לؚ__^�P�MS�d����KIN����1�;��
�uǂ���:�t�!uv�����*
+��)2%�n�%�e�M����]���I!��=��)�M��/��}�!d��v;�dЯ�M=j��� �l+m���-,�ix�^n��C����`�i������ٲ���y�T���� ġ
T	v ��)���pgd�\ͥ�p�aɎR 	�5��'�?��x g}�D�~�?�3�_&��J���S�s)��^�OD�b�=9a��{������Eq�t�4�?��7.sǂ��u��mCY	t}	�p̏�>���9V<6}�r�EK��H!6��	8����<j�/4l[��4�h%����E���?5o9)^���g����_<�? uk�Q����	�
 4��P|���j[�dR��z���O�|�"���I��Zfo�6�ܸ�;�D��5�|6Rj)?���O;��+�<%2����)7[��Fe/�c\+�E�[9#`z��%�$ʄ<����wh��Y��m�O�\��$�Q��bN��ƴNm�3��e�m΍xod�H��?�5^��[@�WHX2��&��n�W'O�!ӂ�pzsLz���A�:z&����q_?g�5��ú��T5���K�5� !�sY��Jh�Ч<{t��q-����%~BXe��y�{3`A&���'�_��y�&��E|>p7��kl!�ֳ96�X��YY�װ�:�-&J��_��X�J<�柱'����<��4�+?�n���r�����u.�����8�o�#v/;���>�Jl�� (��M1����s������]���`!������a#��јv6�=t��*�4|�o�]+�+�m|��6��K$O�M�zy�;������.�J��=�S�V�@�)�^L�*C�r��+P�]�Z�UUZRh3ٮf�!���nFMM���B>�_��T��j�	�jv��_���mE������k�-f�/8r��9�ŋ}Qj�>����N�_=iԑ�$Х2��9�mGr��a!�ط��Uh���^�zBMW��t� ~4/��&��{,T�'�Iapz)��pw�%W��J}KP)�0�x^_8�'������o}�5�ZWq�ŏ�l�x�(�q�QN�6ٖ�)ju�T�M"mZ#^
�~늽��a] Rߚ�u�c�|���h�:�������Z�)T�G}Yr�Xջ��(�)��f�s��C+��_m_rw�@ٓj8��`����Kw��v*~����w��7i���ѣeט��W:dD��&�&�Hޭ�Y>� ��++30�읦%6��Q�}��dٝ?�.�)ӄ��|��8��u����`� =WYP�$.㰳ٴA�R�X14<�6i5�[���.��)�h"43�U�np�V�d�"��¦lOj
kL���p�I����"��������/�uW�u�+���A�H�����O>���]�ػ��y��P��M�N��:��G W<2n]�^���O0 ��ۑ|ʤ�d:�*�Fb�t}������A�9��&���J���$��ځ��ܽ����&
��p4�Ŀ x��Ťx!�*"h�r"�Q��ݴ�����Q�苚uv���r�4�ZI���	:9J�R�L~�՘(��T�r/a����ء�Z�4}��C��V3���n�ߨ�"/�Tڃ٫C��B(�:*Ȁ&�j�4˨����Bl��=m�_�r�?o-t�R3�I���HP%&ZD?��?V%���)�=�uXسd�'����'F��%���t[@��RIVǪ^ʢ�sQ�*+8Y�e��Gqe^|p�'�dDzi�E��:�ey�#�UgM�>�B�t{��}�:�2rL߫g�oqfW&2b���J�g�
U�q6Zu���/U��d��B��f}��U�X%Đ�i�r�=��S�Po���-�^9o�/�Q�|�$��$���rw�8��<�-t��ւ���S�a�l�R�eg�/��=�,�����������Yo���"�+a�|�'q�)����'�.����d0On�J�텑�^ &B��j��zL�X��p?�I)�҇��+��Y�g�G��x�+W�^������ �5p' 
�/w�b!f��b��0f*��ϥ���A�H�q�� 	>T�e�
� 8�2.�s��1Ç<}O٬�+�^ڒ�uM��4�c��7.��N �m"��fG^A��dYDd��C$�zT��ݶ��ji����܁� W�G�����~�"J�{��h�	�D���v�ٽ����!����}+�,N�W�d�Hт,�X�v�c���[��G�P�jY�b]L�8�D3ִ `��<��a"�c��;a�n�u��-3y��T�}s�1��s�b����n�v�
uջ�#�p�~����������}��F��e��-|(�W�J���8�\Vrt�cr"儬�Z���B�o�L*���2����J�=Ǎ
D7c� �.A�O�=�9�:������������F��^��L&�~�MB��ueΝ�������E~��^���'��p�E�щ�Z��Q��'��ԤVU��콾��A7Y-�}WY0��#5�!��s��\��*
�Kb5��x��U�{_Ce�5��+T��w�$ۆ^�v�v,#�ߺ�������5Jr"\x�h�BT����Tv��s�i�����*���1��Y�MN�Y�*��gG畋�"�ʉG\1����?rn\e��"Ha���{�����
���E2z��a=>��w'���'d��gJ�e�!��R!�d�Z�C��F"��&ޖ�56�S�du~z��e:����Ӡ(UZȎ�)��Yp{{��
XQ٩���^�p���`�>ފ#K��_F��5Mr����~B������$�@��! �@���y�c%�n$�
���:	�doݼ��d��<ÙۙJ�H�g���CVV�����@�-<'��-Y#pM�ۿk��r!O/�K�J����e,��^.58��NZh��I~	�1��{�
��U%cf�<0��Q�~K�H���Dl��J\]�3Σ�3�\ئ�dپ�,�Ӧ�6��z�^�r8K��X!5�m?ft��K� AΙc�*+]�#@Ct����u�3�©/���4�FT-��`�ȑs���{e�#�ME������G����iܲҁ��U���e��-�33E� r�"b�|�G��2{|��[�=��SOµnv0��pe��C���]$p*}5�D�?���eS޼��ܾ��Y��#u��m���xv$�DQ����oث@ImkS=���k�"=K�j
\��`-%Hc�?7d�;�p�F��	�ꯞݴ-���b�B�J��W�!?�JLUt��zo�/�=�F���t�G�o���㧋��-@�P���?#��A����0�EO���F�6Q�� $������\\��O���E_)�6�h� ��w> �^��t��n���M:@4�LϘ����	@#�}c.�p+�	�&��୐�N^�#�����V���:�ʳ����V勋��� ��H���&!�yu)�.FdԸ�E���־����U;��Un~y���K��1uRlX�e�ᬌ�Q	W���Z}��n�@�S���{�QF��m�Y��I�����Y�n��w�O��aJ�vfZ��R�E6O�	_Ɯ�Z�^���tgLY�>��o8��nqG�y�E��ꜛA�`����g��W��V�'�+��� X�ϵ���+�l�T��I�F����v{�Se�}���ߩ|s�H#@��|V;M�^`�Or�*%��� �P�Ce��ϳj��|�Ŀ΋����@\u�N��{�	/��;5ԋ_e�<��2/Я٬/!����\��ٙk����sKϮ���2���tI��f��Kc�A�ۘ|�Օdx�"C���5�(���Ag�����4MI,M1����NH����C�6pF�� �w?��R��^AZ� ��!P���'�x�����]�c�ieA��kD"���!0���S��[�������V�c�� �������E6�l���n�������Hv�5��S6!�	a��T��&]$T3��ْ���F��=+��xE���h�H�TY��L�ƫ����3b�u0X�\�4�U�9 �����-�����:�;�5��A8($̼W�I>�8�М��Gzݨ^F��xwE�Ф|����r��>d�ss������
o?� �_��\�#cm�7���<�Ui��u� @<Rv܊WA)>���O�J��W�D{V_�C�ݬ��(Lu���
�PT(i
됹�6dULef]`�lӈrY��Ǐ����WB�/��6�j�Ozl�4��UTp!å
A�5��2��`�a�ͅ�h]L�MO�?����1KD�L�$���e�@�p��Yi{��A	���s'�A�,�էQǫ3���K�����ߚ��ۣ�أ�4B{�y��5+UR1�X9h�~�=��B�e����d�-Qm�����s��>�o�I��(hcLjgcC���	P��gс���cmd�w�-�%�;R��V�$��3���Dq��Х]՘��I�hB%K��C)�����<9�o�츍�˃y��g����~z~��v��&��3�}o:�&��'Mj��8�%|���J�ӑ��L!�D�0`��h�c�d����v��N��Iw�8�N(�%P�r��q%�u�����t���n�p��4�t@��&
����$&��S�vp�\���6��+��(k�֖M��-~Mh�|�P��!(�G���Q��Uw>Mp��wC>������,A0m�MM)Q��X#�n���5B@k9�њz��񧛞-��"7�%v�ŕKm�w�� �B#�`]�{��
�]�[lJ���VU�'�bw J��e�؅�}C�u����a��������ig����gZ��<Y�t q
de�V}�X�@ʧ� P���Jl��ܾ@_a������Z����2�L�)9|�@�H�m�W����o�l�>�A*�z�Rz�M@6��c��x��v�Cr�q�/���zly��ݟ�[DւM~���:��T��a�,TP�?3�����n�V���3VQ!�2�$*az�|{b���k�罟V��^��e=��˅0My���]�>dlkE���#d%������Ps1�l���ai��S/	�A퓳��ol�w]!Ƕh��-�ĴA�u(�
&&�X�a�ΦJ����+�D�EJrK ��5�T���_Ⱦ�w虀g���'~<J[ٔ�m���`T�mΘ@�U�J�q�ٰN��j�6�B+���c`a�1t��sw2�,:����1�_��u�Kd��J8�b3_4^�ؔ8�!N�`~u�7�Ͽ���
��jnJ�	���6aB��;�`�K���'j��L�#ϭ|J~��ϓXoˮ���S�g��&�E+^��I���[�-��W���)�V�ML@)�I$UK�i�d����I�䐤�f�@��Q�
3#�q����9v"�W�-�e�oDغ�|��7+��@��C;�rjh�&|�����2���7Ä��K��rN:MZL��Б����[Wp����l���{�U��u|.f��+Ț���z�m�S�'�*?ye��9&pꭹ�e�I��%�3�P,���/e%%��tr�+�"��r,��u��Lz�y���g����T���P;c�d�&ȉ2�����sa�P�
7�&2hEg�I����.��s>����'��BF��A��d�q�#��Y>��(��6-_�	��p�(��&s�X-�W����&7+��X2]ɍ�L;��[P�MЧ�]�y�]̵�B�����k4��鯙D�pS�M��M�� Z�r�~t� �d�,���Ww4������W����I�,�/��[�	�-�F�G���}�'e�!���'yM�~��K�N�yL��t�L��T�CVko��~�k�����]�	r�g�0�����R��zV�N��Y��7�!A<s�9�11�݊yX�[-nJ�o�D�,�E��ta71�н-��!�_���K��F]g���8~T�D�-�IA�aj�)_CfwO���귻j~�BP�_�?�`i�=l���
�֌�������ܴ׫٠��a�/�y�8����(�QUL�j_p�JK�F���x���"��0��
,:�������xw��d�n���ܞ�Ϲ����D�Jj�ژ`��lb��:����}�Uz�"e�P�)��b���K1ö�<�W�Xh���=FR5������r�ܳ����5"��<$�@�qo����$au��C�>ڦ�CX�����-�çDy����{Ko� ��k
�%��,`��@�ly��j��v;��dOK�Z�Y��5ە{]V�&�*��֭��+ԭ�7� �{һ�3V�w��I�;f줍?�+��dZ�E��Q��¬T�!�D]3�)\�3�B�d�F���m���Es���q�wVO��E�[����%f�ͱ����?�qx;%C��
��0�(�#���AW���?T>�_�#YD;�j�Xfc�P��BFז���D;I2�v����}�B��|P�@�a��I7���R8��α0>|p�GԚNr<����g�zR`Wq��9	"Ӟ�+�	����R�\E3���ME��l7a�+AE�~×�e{��͜y�*�7�;O�}-K/�B�~b���mi��kF��㾝��o�-��M��n˕Œӓ���jϓ�'��y{��G)t>�IE�����	-$��3��}���<���Ҿ#.u�c���ڝ�kP(I̑��y�v��n���[nJ�&,r��qQ�3�:�BC��J���+	W)�K^�8��G#?��h�~�Ƣ��3���|d���K���V��8=�1�ǦG@�p�S�oN�����8M�f�?��f��lx��\��zT����W��]l:�	�]B"2�%�{����߾���2N����S�����q�|~�kV�ɺ�-�0y���:�<�g噻����K/��I�M�uaG}�_��S͂����ܫG�������[�bE�n��k���a?��(�q|���Gj�P������)�$��3_E�7
c%]Nf*�ϵ��wH5- �_mo�b�U�2��7Dۮ�U��|�$2>�΄OS���Ą&�.^�����x���*�z�Jͯ��>��ɚW��HW��<N3���j�l�dѸL���0B#ۖ*$�ʃJ��.��j�%�Sz�,W�c
8\Lc������'?7U�d�I�����N$U������δ<
ϛ8/���%��G'm%!�]��U��*�1�d_�~�V� ���	A予[�؏+���˴|�asr�2�S/�������lY���.�Т��K�{��)G���3���c�����
�<��3��3��@(�|��d�r�L���N���M��:B9�~ҫ��4`~��Z��	A�X�����e�.px�<j=@+����w���:�NOhn�GOH��-��lHxV2�=�V�xeO!`$7C�b�z�h�X�Bk�m1s�<#��T7g�E\d�t|��#R6;�������P�w.�)e�T��q����*$ s%)�,�n�|@�g*���`>O%骘k�f��[��~��� ��P��
�����,W�[m!="	��I�/�^]��7���T�Q8�KL�^R�V-|$͟ȯR��n�[(��8۴���q�e�C
��e��U�K+(���o�:����E6(��Ǆ�j��<���Y��	�c��)��6�H�p5�cѪ�V��#�uc���M?�l���<?-��b`~��ө��7#�v��F�ňS1����f������>��-�Θ�>�Ԓ���h���ݪ�ڒo��2e0�mb������.���Ӭ���+���{w��EP��i�HM��`�6+{S�����7�	2��e�L�4��i��f!?�h��J���EQZO�~�M���߀=S��z�SK�zn��H�F�x�-��sƍ'�Og�3�|��R�Gcۘ׿l[��W�/��Xj���n�c��=��c!�,�r�h����R�jJ��HNb��%to��5t�rEc�v�vO��9,��Ȥn�D�^� ��l�M�'��yJ��G�O�q?�{��"�X��Yn� ,��'��GA�#�������`Nۃ8��T��A3�[:���Gl�:V��ڢ���ک�5��@���`{�t3^��]�5h�?zz
�k0(���4���,�W]&mq���h�1�:��q��i��M�����;D&�o ߱�.��*v��c�0q8�w����bq�����V�KLc�Y��o�4Ks:��Rd\�'=ߚ��Å)hOFɩ��ʨ��';��N�S�<s/6�hSY<.F��5\�sA��o�9j��kc$��ՠr�u4��߈j���j��z�)W����Mj6��*^�WO��� ��Z'�!��8Cv8&v���2BlKk�j�Q�1��l9܎5>2	�:��(c~�J��I�>��>��h��@$�qkA���ŗ�!��uD_o6~8��VO.*@#�YKH���>�s�aV��
��+��F{�p��Q�[(�����]�C�@��z��ĺ�]�(v�oRW�Q�mɅz���bH��;>�W&Ҫ��Ѝ&����T��}��"����Wv���6��=�Rƌ�&�����Q/� uڛ�:�C�QD����Q!�'KbO�qP����L`�U�"jPC�s�)M�g	��v���(�����1��=�bN��͇�+?aJ��҆j�)���'ʲ-�����\z�������[����]9��o�%+��T�_#���Z��O�<F��
���H��RFE];�ۖ%v!+Mj��e�a�i���xB�0�Л��XX�D�{�8�ﺨ'���A��n)n��&*�a]=���|Q\V�޹��^��z�P��qd��l�{����՗L�]�ۋ~��25�jbr��cZ)<�X��z@�@17��n )��K�F��(���x�@���e�᰻��p�`{tz�bE��^X;j��my�?�0�e\'k�h2�qz����5�"�8�o�E�XlxVHYEB    2039     9c0�0�m�Ӽ���5��;W�|r?�<���.R�H_Uf��N���ٝRQ���&�5:!��?���W�Ʉ0-��=�W��JxAx��.�9�/�a�b˖d�Rz�%�)f)7�P�� ��a�Q'�.+����M���ZJ��	�j�������YjM��\�D�+&�+��2&6	���4��CO6NV�+���.��Ծ,C'���
>�ʻ������Y&�惬�����9�3<�vW2�������BV�����niƎ���Hn�^z[�lR�lp&�?Ն�B P��8yz���٠t�ʿFW��C6푖�����	�>�$:�WG�J֏(���b�.�;8Mt�m0�c�����M��Feǉ���"z�����a=\Pr_6��!+[X�U��w"L�M��@u߱��f��l��˃���.��*�6�9�=g9~=Y��J/����»1
H�nc�j��R]�C����J���/�{�����m����8
�����kJ�m�ߒ,=a	P�J��g�F�g�����;�&!���ثŬ�|h���^�gg�4S٦y��q 5������B�~���g'�b�!��W"e�Bc_nԚ��될�j<$͉Ec���I��x�S�'��Rg,0���h$u5dz�~
��~� s�!��s��	9���gE?eГ�<Ȃ�L�v�P����-Ů������6O7��v�F+���=�^����`N�=`I�R���`��'%*!!nʁ���FU�u7o+��KKĆ�
�Y�^��,�S�C�� B2��D(�D�EC�S9�{ˈ�߶n�lh�Q��>(�A��M��tx
�B&��G9� 1/mӗ2
wA/��[O;Ӗ�<��`�\�aY_��~S�����+�@�
��h<(�a���|����I�a4#d(k1�G�ƚ��:���DW� Q��Kq��Ƭ{�J��c4T.�x��(��]�߂5�J>-U�\T���7�15h��G�B~�4�pFeK�霘���[�Rߕ7�p�qȓū��D)����V��	�C��y���)���#õɨ����.G;7#c 'A�<��( �3s�yq�d���k��U��B6`J�q&r*��>%���ή��:��Q����<BX4��k3U�3��Z-��Z S �f@ r/١�K�%+��pj�'ή�*|z&a䌷�ͪ�|.PB>��P��M��>�HY�!�fe�HBl�3N�C����]7Dޏ	�^t���ٜ�7A���Z���Gq��	��s	�V�s�<e����M/s���1��'U�ZZO���J��=����Sm+�6	�
�jp�K�L�[�(� I[�3���
H9�'���ķL�T��㗇`��J�K�S̲�L������ ��e޿莛��_u5�K��jW:hPʱ�.7���!t�K.A
�@�ޘ��K�f��x+c�J�,�шb�ej$`!�����e?�=[��^�����p���@����2G���h����ޱ�p�EH�~���%m7������U7*%w�i"h���)%q-�e����Ҳ)#�4��h�"x�G`Qу�������}*tҦG�܁������kG؅���,�ӻ�XZ����^����:���9!�0�^w�c���N!zL��ŅYp,Y�4�Z�x칋�w�.Fb�b.�9���.�YT�߂��i;E`�ĘQ�V����Y��{�yHͮ�S�bc���H�H�����&B�&O�k�A������/�&����z�JQ�V{n�oBD7-O�|�	��4�13���֜�c�{*׍�u�2e��O\���D}� j%ڥ� �������5��2�f�Ku�)Y���ZH�(��*ؤ�z{:��و��Cx�t��0�	|���eS
O�`��˨�1k��!��˖�ZǞ��ﴈ>�W�4��\�c"�\��K\���g���w�kVLo,B-�������ڀ��"��J�Uf�e}V�`��5��*׈��=�L��х��BԊ�	'��H(��r`�d���q��r�:ņt'�����j�<P���"�ܔ	�<�C9�'�"�&V�M�*��n�Җ%���[,�˞Q�dfa����K&��P�+�%�3/_i�B핦�m��@f��*Y�0)���Ace�Z��v>J��"]VQ�[��U��>��o���3�"��3�8xx�	s�<��S��.�y} ��O�m\�O-��S�knL��	�y��E�۹U�%v�v!��'4�9�"�7���B��2�US�d�O�x�f����]zR���D�*�D��Y{��F�������A^㳢�Y`mk��C{9/� ��̂���-c���0�F��-��>_��E�`9&��*�h����f<0{���ؾ\n4i�"�m�B�"�93Z�H4·�ԋ�8q��Bj�'SW}�ߝ���SV���v�>���	�O��hh>T�]p�