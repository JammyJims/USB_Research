XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Vx��p�e��o��y�tp�M	�W��oe���I�8]�G;ܭ�ޣ�x��F�zCj��FͰ�)ߠg����q��b�.|b�Z�����P9��%~�T�	ז@$L^�o��Mh�7)T����'����{~c��j����Ȧ_����
�e �W�^�B@M�_!��V���\Qv �����8�=�ru��i8�����:b � c ����4X:y1BbW����.2�~�B3��<����H��1�_�v��3������k7�׿Um��]����%Љy��!bu`�!���s'-�|q����
j[��,;/�q����,u�ffɌޅe��g�KDt���!����#-�^��Zw���8p�Z�o�g��-�BѤ���k�pCQ߲�)[����D
�NW��@����D3aw���f�0dJ9�-\(
�����]��'���
%��,�aj���]V�~�5~��)����gT	芏}�޶C�F�3j-v�,\�hjz5�35� ���j�u{=9�c¦ձP���q��	z�A�,�̱Ȑ���Y��1C�:�|yYQ�����S2k���]7}�
����������%�]�y��	�W��+Po�2����x8]9P~�G2�j,��lf�6�ߝ�A�yvYE��Y�V=�xv&���q?%�J�[IUv��P�o��.�)B4��E*�V<h�h�%�Of���\�Rk=��Sv ��OiDE)	�m6���d��$E�
� @`��Rl\��XlxVHYEB    559b    1100=q@�P2;�R�����\i�&����x���]F$���G�tX��ɱ F�g���@�����O�m�x�~N2E���t��W뵘�n��x!(�=�xp'HqG{�,֏"Q0M��a���������͔J7�?���D�o���5��c$�5g�~���{��{!].?��Cc��<�>�
���5
U��(��	k���1��|yM������Y=M�0zR��#�A�LR�e_��˧!�qo��>c*^n����D�l$]�Q\8����Gx}�O�ČBE���8�^�*�Ǟ�qc��N��#s���N�cG:�'ep>�T����;՗H[Ӷ4k�u� ��k�o(s�\{J� ;��&X�����{-����������1���Nk����P1E}ե���m�Rn�c-�l�q�o���<x��_�&&�9�E�,�)S���=_ɩ0��!�̲-$�!��Ȑ���l���{!��A�����3g�&cvL��"�M����*��5˴X�k�ϵ����s�ڬ��ޖ�];t���H�/�ٳ����k���h_-�<0�&伝�/�L�9�]o���'�汇�}x,d�[�� Bj�_�;A�+�Aƺ��{Ns)��߾�sgNt�_;��\>�.E��B�6t�W����j@I�4�����G0��<�-{��g��S+O���1V�Cv���y�T(�w�G�岓�u�@U����+g��N��&�����~7g�2��"ҝ�<)��e]p�wоA�}UDZn�ݛ��1�{�{IA�Э>�<�˶g��MV<ӭ^��	ry�mu�M�J��=�l��u�����Ƥg��6��(�X� �Xm>����bҔ����)��n���D}�d��i�~�ƪ�y��BB�?̋#�nk	��DFh�Y��Y'�ܸ�?�I�<<�bײ�+��P��'�Zl�Ŕ,`��Sѽv�����S,��a�h�k�ܰד�[�+O�`�O���J,��ZyS)փ�xV���LW�xfS{a~��HjD���7'Ya���0��y��0��Se�7�I��}1�1/��W�M� "zك�4�Fe�w��n�����ϐ�k���X7�m���+�{�,�+40*���\^��
�U�������@��{n��2��{��b�@�r�]���C.)_�rjޗ	�<����L�v;h���B�S%������a��J�r�lp��_c�a�w挣�_/R�O����L���&O������[�"��D'���l��]��m��㶵�H�T��G_���q9����Ј�"��ᅺ�S�➦�\k�K�>���y�{�:�O���[L��O�~��|���Hٞ���I����c��#���q_��ʩJ����4�\��+f����	��K_�[�|�N��>{;zҕ�#�9NHs���/Ab��g(�����^�G��˭��v �;B�c-�+���Ƞfi1��V���C�-K�-��\p�V�4���� ^�YF��m +X��Y8����(��0��#&$o����WǼ��q���Ƌ�f��pkB$i�VU�LsM@�V���74oͭ2����W�;/��QzB��bJ�p[������0�7�
03� /��j9��?�O�h�}5��%�ۺ>9y����a DM���\U�+���~=Eiw�o;w����mOխd�>6Z1r��Zw�&�_��/'��F�2%�e;�[�E�Ҿ>��&��AhkEw�B}���ns5�w\9�=�jѭ���}VTP&�@�]�v� � �t�/Վ�C�C�.�?��CQ�h��.J�[N 9���)�|���/�J5z�k�^@�8�.e�?z��#�G~�tw[a!����9��݂�SJ�@����Lh΁�F6�.5-@eK`,t���pp�f��$�y�z��<���Ӹ�T���3?�eť(Tpk�V�����}��k�����۴��?�!�O�oW�d���oakM���oe
}�=$W���H�W%��ԧ��*��;�a4�:	��#T^�q�1IT��B�v��⏧Y��X�E�Ap�;T��d2Y�g�yy�6܌���k��q|�8/b�������O+9Έ�{�a�h��P��o�{5V�|W���U8�	���x`ZK#�	I��eU���5'��iL\����VW��|��:_��M:XTo!<$����iI9�ר"����p��Ž� '�x��@a����J�rv�x�PCc�K���(Hр��"W�f���%��B�c�^��GF��������=<ǔ�:I��M�qo��Y{]��Wv=x7q/�F)�`=��4yTI���:�����\�������:at͔�k�ѵ���$%��6�����:aB+aw�Iz�Q���`��f��Z�TU�k�z���9id������ԌE��j��}:N��W鞌����y�p_�������`KU���k+�1zN1�(b�R\���{+��6DQ#�G�r� �#R��:t�G���o�����?���8?KẌ����Z��G�|��I������-�aǹ��׃⼁V���mX��ܮ��VuP)���6̐C�ޠ��ݖ�ld�!E?�����Ž�%�!B�}��lGh�����}�^%�4<�3������� ��#��G��I�W�ݷ,@oR@L
D����J�Mq���sC���I����d��F����W=��~�(���	Ay�i\�D�<���j�9QfE���?M��� �m�a�O�%��tL'�p٤�[U��� aJ�?�I�]çN�d.^1F��IUW�8�k��>�+g�z��^-���%��/��뮿S󆽉�*�O�dZ{����7���,m����_���O�V�<��$䔣m�H7�]A%6m�+gI��g}|�u��kz����Y���<�O����M�R�h������`�t)��2凭��5��1�{�q�:K�8��w�%q��ղ��ՒK�8�-�e�wߐ�	�[o�T�����0�.�W]�&6"<M�Q���~ ox[�&�Ds�r����XO����a8��!��t���Zh2�z��
V����P��6V��4�eW��T`�A��瞫�:ٲ�~p%�N�0R`�UO��W'�I&���:�#N-��wF,������n�<��I[c�ln��],\C������d�t~!�~�[�ǒ�����Py�ͻ5a�L&={�_3���4C�O�����2�P�9cS���&%�68����YTc��lteR
��|�n��EJ>��v�UJ�e�d���s��W�0�
���猤�E�
9/Oj2���q*��Y�г���}`3M�e�ɡ2��*��1u
�B�
c0E�Ґ���%Hn���/�yZ��.���ʌQ�-�¢R�A*��Ʊ�����Н&	O��AP�D����o������]�=C��<����UToT;㭄~|u�(���E����A�gR��X��Z����m/0$�56zW�6�Ƹ��v9�;��!eg?��-��]K�]��&+�m�u"�B�`���g���K�����[�^�c_��j�0n3�a�8�iU�Lb5�7b�^�T3c���
��������?񃑺�#�7��Tl�S�G���hRue�'���4�f)7�$�@/h0�L�1C��V��Q�܆�΀�'�b_��'�68��_����M!�q����`�1��B�\�
'e �\�˔6#�E��s9pK�w���>]�p�����ϋ�����(�}�M�e�#~�����=n�6rrΉ��O�f��<��9�z>����G�4c�*���� �&x?�gŠD����_�釶<z��n�W�MV�u:���']�3�c�zq5���^���<�tP�2r�Yqd`����)��Ӎ�.-=Z�wH���E�e����b��7��ūy+5UUq-֛n]߷�WȿxY���C��>���l��cC�e,�y&���'�k��g�=�����	C'�Gk�S��N���&%��h�u/5�3�
�2�ve�����;0��N.v���>��@�p��d�����ϋ�r�A���TUb�ɤH|�f���e�������$��# m[�T9E��c������U �[L�-v��g�A|��w������69���t�����\�AO�>��,V��$�##�3MFD�I����e>$�&X��f򍌍�a�S�1t]���0̺2O��<Y�� �ȬJ�a]�����B�t�4�?��R��29I���D�C���PR��� ��D�FG���k7gg:������7\����c��pea�