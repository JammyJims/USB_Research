XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�.���mh\ƫW�ܬ����򪂆���!	����=M6U�9o:�!�h �:.�K�.l=Hk��9�淰d'f#)��Ú���,�V�G�.������S��ؑ a�,93���؉*��_GD��Q��!����F�C���4��n�m�p'�����]���ҨW�����F���ľ@�dP��}4S�d�Q�Q$��?����>����h@gE��*֡Z�A\y�IAfJEs�!Ήk+:t�YN]���>f����MTϢ��D*��(O���ԃ<�������y��\y�({ԡ�䣎;F�=;��{C� x�F��HѼFF����pII$�񀁦9�3k�my"�����E��ꅦ���_��c�c���{4r ԕ5��d�1h��OL��I1������ ��X��I{B`���F_5�͠�d�VsҢ���ޏo��	Vkt�Z�f�)��*7�ɛ��)��ܸ�Sɫ�LF�l�f}Y�9�F&�KC�㮜VR{�	M�贈�i�Luv�f�t��p�t�Xǋb,��&@��f���^�����]�H�H�[�(mf��	�R�=��d��LrB���*P���2{8�<�0�2z'+=񯰏�!��Ps�S/��J�Y�s>�0_�z�	r�=?K�)�\����,���nO�.c�*Jr�΀tJ�@?dA�*ڨd��g��҇/�o��{�:���X���D��7��bj�=k<��:�	,��2x��}+�/�ƕ	'r�BXlxVHYEB    fa00    2080W�ڸI�B�F��.(5��4pt��c��N-�"�������K�][�@�����s��e��fW��(^!v�L�飙[����H"�?w$��e0{�=e�@{�
E���Y��B�:
��dJ����!؍^�*{`<�H��0��ei<��쨷qK\9���� ������
���Q^�tFC���א����=SV�sus٣\��j�8�[�=Uv"*��cj_oʚ%.'W(l�\{�>k,��d��9��,�*��v�Sl���M3�7�R�=���X���)��=[�t��B	�r��9!(�)(*��c�F7�ıe���(���j;��B���h5��̆�����\��i�+X�(�E�?��S�4��)q�aU���ц����xVn����jt�<��i�MR��K����蓸�f����۪CW<V�����5r���Y'd�ks�/(�	ٳ��}�5��|�~�*����{bvPp7��Bm�'L\9/�cˆ���D�y��j�oV��r�oU�p����2��~�y¡���,U���m�Y�b�~�iVcQ��;��T�����+�h�0�&���� ����`"���O��_�MyX���\�e��b��ƶ����?�+YhI�p�֛����$TS��<���%���QS�΂;����Ld�������?+ �c�]�ᰵ�J>���w��?d��J�|��sJ�h��D,K[J�U�+��P���r<���v*;��l�V{؇Kĭ�ۆ��!��^�&���ʞ܈#�ڄeT���|rϺ�#�C�?:�)�GV�	;���J���D�~�g*M.J��v����l�!{Џ�����&�.����K��"�#<���r�E��C#vͤ�����V�����o>�e��� ��j^����E���VE��'���=�i�yaY�~]�`�[z���g��O:M��*6���up��i&�w��[�hن�U���]o��u�"98���������� ��;�ۘ�Q�ʹ8QA@�@���b,f��{	+��7�vg]i0x��/ib��Z*���9��By:	��WY1���j� �.�N���&�x������~WY�Q����t)�zj�������$��(wjh��1�4v����?ir��� �ҿF��K���ʽ��^Jΐ�*�!P��*��B�4�[�-�8�
�,�f�H�)&\Y�4&��@=L��X0�|j^z>�洼.�i����b"�[O&��Z-3�_��~6��
?�-�Miv�;�i�����$��s1��%b�e+o�'�0N��:' ]�(�2��/�V�H�&�٢ވ�3����{�nr���K�_0פw�5���^o����+W4��/؅�c'j����NM{��F��U�-]3�c1�_�b��˒E۽�5�RP�m -)H�U��\;���t��<ҝ��v6�b�)A��R����2�x�A���HV���G��t�8[�׫}��x�J�%y`�J-;q;�TF���`8���(��`E��ju+�ݓS_)��HS,2�~�\�|�5��iJ��$�9a�J2`T)]J�2�×DpD��1����X�o ��C��VuDd@KO$_$e܋����=�	��
����ou�W-�/�k:�<�ӣ�����l�����]���<(N,�v�&Q��w��C`�re���ʚ�e�A�i�"�H��HTy�>�#U�2;p>��3����`0�D�f�pȳ˔��v���(���n���Y�P����X��L�b�����P�@M�܌��aq�_M��I?���գ+l�b��I� ����EW 2��Pz���6�a9����*�	U�օ��㢜GԺf:���~��xn�lm��㑦Xn��i�9s�RE��\nM<�-����9��V��Q�j�s�+���T��5	��|"���K��
���&�P�>8(G1�&�٨ ��1h�5h܅\�]pZ��W�z\�}����)P�1m�5�G=���v[/a�y�7�������7>>3�i���������t�~ _1R�P�U���r��F�a��˧��-��sN"x��Oudn��L�u#m\b���O�D. ��e|����nY��K�����{�f-/K�O[�h/���2��фA]�1 ���X��V���^�Ɵc<%2�Hi�}�o�)�҄�9���(�X�)]-Ǭ�ź� 1�i7�qFkz���ݚ���8��5
w�U	��(�<�q\�X�0���}X���a����J��2�|�@.�[� �o_]��w���8� �u�x�u�G��0�q�R(��Ymŵ�rn|a��8R��a+y�V�R_� ��'����7Q���SldY�ū��i<MKe| �pU�%�#�~#�Ė��uֱ �Q��W������,)�,:~��R�	����V,ݱ�2,��bd9WWr<ȥ�� ��d�F)�Ud���w�S��1�ە�4��1>!lK3�.l�Ʊ!|��!��ϝ���/�������U�V_V�
���2�t�n�L)���&X�҆��e��� s�c�1F"��j9kG5�)<���$<Y�ۓ%q�o5m5��*�id％bg��jx�x2n�ܱ�-Z솱�m��󥆏��j�����lh�?�BH��p+���l�/�ŕ�1U�\ jk=�{��Y���ص�1�Q=���D��1�D�4u�W�À����@#{%-�p0Җy-�V[��k��x��
��as.'����=(�2��J{q0���J�	�����v�륳bGH���$�I��c[��4��C�$ZƲ ^I��9Lc�l��bZRq�紙�wȪN�ĥ��}҉�n�i�Zߍ+��H�躗�f�K��>���Gp�'m+���X���0j˽R` �Vo�GC�ᷢ)9_�ĩ݉x�ђ�?hv�港Z���&(+�h�Y��(PK�=&q���'Q�18f-��_��������:8��Yt��=���JUl>g�� �i�Y���OI{r�S;�����wOC�5�{��j����P�<�F��Z�kT<�?��)�Td���[�.W���=�B�K+������U JF9��L�L>m�F��.xq�Ä���)��A�j2)6�[�ʹ���lĢ�}��u��~z�mWb{���&��)s~l��e�~�k\��}�W���[���x�%�=�nB�<��M&b6��� �ռ���K<�:��Ԇ�@7�U�L��ee��/��{��u����e���X���q�����^L��
��H.�@f�,�b��&M��,�@P8����x�5�0d�&Ee˽Y���E�;y��8���Z�	y_Ă;	�����g�Жlb�+��G X�&5�$�7��ʅK����i��3�9���4�Q�J��2Y�n�btx&�"�g��[ԗ�S���i�3*A]ݒ��IMF�����Af�Z����n�<�	��}m&|����,ë��gR�M=y{���,�'93X����Λ�Wq80�sa�Fm�BL����������d��%��`��l��-j�����9�(׌�0���Zj��o�:ڤ��^�����c��D5ѐ9���n�	�M��(X?*�dR�E�����=����^��دZ� ��x�}kL��L��w���W�����"��������LwC=�C�د/�@�"�Q��6�3C�L��,I����VC��?�
7��?B[`P�A~��ϙ��$i/�?�|	�[���4V�y`s?��?�
�>�#/�u\�' 7�Q�7��#��Ol�KE �}W��2z�K�aRv�	����7e��)&��)| z'$HIH�bú-c����1U��o��ʌ�h�qZ��y�������\�sd�4E�y!]߻+���l�[��A�"�BS��qJ�K��R"Ɲ��q���Ef|DY���:f�L=,�k�Fp�H�[�S�gT�����#u��`��Q�TG�P	_��v�̤��- K�n���/��N1j���%(��Xh��4�|����.��U�����22ִ�3��ӻX�'���WH�g�Y
�WJ^�|�w��j�B��u�1�����Fu�S�E鮈�F�O4���Q��E{bѱA�a���w��~}�C!��_1.݁8૱e�N1��2��cV�4�1��Ӗ��n�w�2�� ʦ=4��� �X�H����9�I�Q�s��!B*^�,x>'u�)������,+H����倡�%0fĳ��T1�f�e�	o��418��+l����.�.�'���w�h�OQc�V�D����9X��_%Pa9z��ǇynX�����!$��oW%���=1�z��Ka!�P����N򡐦���8�aJ}4�2?�ͯ��2�#�^���w�/_�@�/����n�9Έ��]�$��J�����!��+a���pp�@�=?����P�W�o��Ȟ��_}j�$�~���ā�w�����bR�rR^�GL�ۈ>��m��U 0�+-E�U<J��9���Q�E짵#N��划i�-쌗�)�ت�����~lǶ�8�[�ү�%�����K���+B�;�o'=��wg��w?1J��ww4�G��Ew���1�1��J ���U��K�5B�̧�B��A��J��/92�f��W�)�~<W�1��5�X��[�	����g���1�R��r~Ё�x��� �ˏ؅ٺ���h$���w@z�H3�3�`�2�>�Y����ma��y�ə+�r�V4���az(�t��
ĳ�?������;/�S�`;��=�s7��z,�l<Ѽ6pzf<E}�e@'��p���F�|�(���B�������#a�r��c��Le$,be�g�Z$�	�ԥ��4�$���1	;^�5$�;r��������t�g���$|��h��$4U?�ba��q4P��9��x�{~�[O��g��T^�b�[�R�}�~p� �
"*֟��s���h����T�^�Vj�?'��X��̈�_lh�i�N	]Õ#�����	�KqǙP�:@/3��i�Qw�Fvm��]?jҎcAe�g�%f����jr48lO䣮^m��W|���,�������Y�{I���[�F��2�]X�(�~}�וC�1c�b�)��8�Vi��e�ts�D`7E�D�q���L���Dl�ae/�Oxn�S��Ů�o5���AXU[���s���O�<��O�!�{��*� <^nK� =��K�pHI���(�(]���2�WHB]�)Ϋ6�Y��K9���Q���{B�ڭ��E�~`�O�71{3ÁҨ�C܌~�t�pz��(�A����PD�D3}m;��.�j�52� �tܟkE 1��uX|��7����\��?U�&���f�$F�:$�Cf���T�]�	�ߓ4 ��BwwZ
�N*Ȧ����aV���i��j��ep�8~� �u�Lf�F�{�q�=�"����Q���u}�z�O+ZAC l�)�/�e���Νz~q��\�
�R��)Y�^��!+���S@ ������H�\b9�Nf�V�i�c�g�oP9�V(Y�m.�\�ORA哠��4[�<��eZJ�ĝ��&J�KKinڵ����@S�1��@V�&`�V����|(�<����[A$^B�*�"�
t�߬��6�/-yR>�|�o���ƻ'#�|m�� �yFr���*��?�N���Y�ݨ�}��j�S�,dx�~?�я�]G*��뱬9�N�9*�9�-���e5��h�/�(��/�hM�� �q��s��1����j�R�t C�W]�o�1a��/Q!�s������x�u�ſ��i��c+�m���� ��O��nGV�a�N�Nݜ@JbJ$���	�Kb̂!�;��B�,��cu[�\ڳ ��H�}�4�p1�� E���jv Dһ �^˗��C�"��n���T�]���H�4��&&.�@�e	 �FA�S�=��7ϕ��'v��G3�{�C2r�RbK�+4�yF05R�Ek�%�)�0���5�ـp�(��
��)Z�e{�'l�t���H�ex?E-�cϩ�=��d:�&?s4k- 侰&����j&�\���#��`��쐒��U+X�C���݌K�?d�ۜ�;�h�{��yL�y��˪���t�<U��$�|���X�Vb(S��0�,�$�h�dge��	�0J6����Jx-�o,]��ܱ�p,�_��t��Ṋ�=/;tɒ����m�r_�ݪ�{[�"k<ܷ��O���*���ő���Z�*R
��p�V�y&��`��̲.�o)��(�!�'	��=um	0ڞY��՗�0�n�W\��y)?@�FGC���Bmu��W�c�6�t5�`�!%͸a{����B��A�K%4�ۓ{(D�_�u#���`��� �
9�z��=K���9�x)�4<�2�n�]�0��	,���ɓ$&
��"oo|���1���|�.�}�pZ�����W!�7�?��뒋|ZY�*[T� Ow#L�ٶ�'�Z�H8 �{?�]t�q���O�Q�?��X
�5w|��o�azX��O#�%{R �/$*Ok���M�W�J���S�q��(-AUk�$��+w�XN$	���Y�]_jR�F7�E�ש�UQ�|����.!�X��ɒD5((d�'XYRd6���$�!�\\�4�7_�ܤ�Q��i��� �P�ts�X� �U\�p��웰����qOA�/���-m�P��F3�o7X��]��D<�C�w�]�����Ӫ�/f��Vu���bL�=MLs����,� t'��ՍkS����[�"���d�Z�G^d��KI�=��9����͞Ƥ{�Q3�v�����u�`B=�T
<>˒bUz.�Ū���Q�	��Q3���/������߉����ċȽ�e���*�K5�'�� �z0x�( �]7�1r�H��.��z�� ��t�Of�/D�`�9Μ�L��r���%9����EBg�P�g���ya[���=���nIK�ޥ ���@�}��@��vt9��!'��b�����31&YPP�HҐnZ9�D��靽P΁����q��(a��i(��}?qR9Y�n��C�䤄��`��Gvԓ��`w�S\j.O��?�B�����ش>��n�;,��$�$�p�� Ș�Cτ[dVx+���}�c�ǂw(}(e?�*'�#��!@�f���b} -q/���촃�o�Ml���IY߆i����t���!&����{)�]����4L��u�K�qRzeӁZD;��P�*��"��Y�I/�ҎYʤ�x�57M�S����cm���G�r���KR�ćgU������=!�6=����u�`�픣V�T�V��>}Uy�� BPt)l{kY��)�^��Cb8��
o�'qo��`_߬�\\�@��"���Y�[b�AHv��W�SЗ�+�r�>^�)5���7��7:�J�3ޠ4�ٷ��[Ċ�`D&����ʴjh�ۇ�����<-)���/�tb���Ӻ�Q۞�Qm�F�p��ȩl�PIv��	�	6#3�R��#��4�(eU��j��	��Cږ����g(8󸺖��ڵ_r�� �n ���qU���BhH4$ӐH[����5>認���	eU�(1����
���D�l��|z����o)������a5���*,ֱs��J�A j0Z�:��������i�j�E	0�ܻ��>Z�F�h&�� G�d�b)c?><Əc��c�d�Ti~ɯ���}�c��Y@fZ+&���n��)��\�����U�����.h�^'<?�L�x�e�Q��U��)���o���VI-	�cs���q�+0ͱ�>����< avؔ� tl��X�ᣙ��*�;�I7��.��,�s�yHiiI%��3��V�b$ �q#�[!���0A-{H�!p��v'\.���n_��@������#��J���B��5���S�_\D%a�:�L���|�e��i#�Pe�`�DJ��T[�r��n��Ty�d��ok��Ia1�[V-��wL���+�ޫ��%C��,�����q���3�id|�j�F}��C�Tӓ�\ ��"��G��� 骫n0�����0+WO�$f����Ҋ
Dm��fJ�1�y��w(��a{������-�>�ܾ����i��R$���5�\�	Z��e�n��U��K`V���]^����F�O��LG��@Osw�^�JJ�֘XlxVHYEB    fa00    1570o��Y��=�̋6��5"�]��<,�|N���(-�˸�!����R�N�ho<uW�=ص�)��~J1s6�@_	UlU�!�@���I��/��Xq	�I��V�����:[C���G�z�b��sV�#18�ϮY!0���0�����~΂�|qg*M�A� �����z�a�m��A+f�bk�;*M��"Ft��+'[{��!/]���E�E=�X@3.�Oq.��xn��5{2����>Q���87���t�U"m��J6�����K�����m�q4�$��ƿ�?H���͆\�1�5�0�t�Z�������{����_H�\_�gP�8f:V���!"�(���!�M]b��vA��K6ڬfV�;��?�
�]�%��t�o�~���*i���<GC�g�����t�fg���l�n����JT7��;�B;�k�}#��q.dZZ���]�fy,�OD(��mh&�a�@��-I�n��a�)��p���=�
MZ�II�2�?�Ċ��3\�(�&�@���4�g�h�QQ۸'����F�1N[��C�5��M��L��丆�\%R��C����F�'�b��$kʒ�5������HH�Ɋ>e8R�P�3g��^����h�sO;���5�b�/�G;1���RS��y����h�K
�%�����|��,4&R�HѯZ��$^��q�w�CMڐ����/ѕ�n�&9b��/nx�J����Ѻ��� � ��w� �s6���{�}l��wd��z���mM�X����\�=�}B惆s=1Y �l��PU��ⶳ
c�yT�u¶k���&b�����2���s\B��b�5�4��9�@+fJ��9���m��Qޘ�FA��#}���{2j����~8B�ɘY�	M��=U//\�Pl�����@��h+r��z�$ܫS9�*(��Ћ�]dզ�g�zч 2N��N:,�� @��y徘g��t�&Wo�K����^�����E�4���Z�Q���'���z�u��̡!�ٲ���b�P 1�7r�n�j���;�q$Lҽ�֦��GF�g�ō"V�W���,��L����H�,�G�B1�g}��_�f�k�4�����o��"%.��~VC��b�=k3l���0�$�ʱ��U��v���
\듢�󘳄(f��J���g�N-xd2mX1�F�P|b� ��B�X��EH�*�U!R�쩚��:���O��~��Z��g�= Nn��O-�U��A����'V|dIZ^j�jtm�B{FDF��}�n �;���3�+���
d�Z��?���I�� +)}V�5N��\V���ffjt�	8f����r͑=(��A!�m}])�X	��1u-z�����t2�o�\���nj|�P?0��:9���F�\{���L*'�_�Qڤ��	�+A��գY��Cr��WyY`�t4���֤z�[6��~�o!?͒�'@������(�BL����+������R�RFъ�iy��>r�v�P����)��15��؍B�T1�����FO�`���8�U��9��5!����t�j�q�s-
���rZ��������
o�EH��;pŜ�� �'F�?w,��$�ȫ8��xXը�R� ��"$[���5go}�M�U��|鎃_�wυc&��[�x���Fͼշܷ�=�a��4	��[� �:m�$[̫o��лo��2�.� �j.+L�> @L�X~G/]�!JiS!�a^����9�pE$zK�
rs+�.J_�f ��Uě:M�ݯ?Ȧa�y�%S'�}g`�.��ߊ&��@�0S�޽�aG]z�IY��<�)�)��c{���u��s�����5�Õ��;:.z �>���W�~�L�ҿ����?vqlL53+磌t$�fʹB��W�zȐ��L$I�̫��M-@D��l���(C���{w F[;$�#����F�	���r��
�<Y�l��k3�$>ވ��
��a[򢴟�=>�r��\3�����4
��;;��E~}&h��Rl�m�A��O�)�I`�G0��?���Q�b)6PKf�T�mx���b��.�-fc�QT	���˒L]"�6�ؑ�����.0
3G=9c 3���D��("��e�xxf�͚�|���FVg�p罛8��s�&,��L���'���u�l����Б30q��1%�h���)��t�2��=@l�tH+��لP-b�ҷ���Թ���!�o�����_��_ۋ|�A�A���XQzޱ^;��9�8�jnX���� ��Ey��� f9���^c�ό>�`|�J?�<�[]a�p�I3�n;�5�b).��R��\6	�������������^��/��>��"�0?�� F�4��{���LZs}�S�Z}Q0�ц��b�P���RF�ݏ!�j��H�W&�g�y���~\�-��wb��^I�3wC���C�K^�F�X�ţ�3.����nk/?�^��n2w��;�a���OF���6�#��ׁ ��J�x!�8���:	A�����g��������j�#9hi�RPF��O���]"�B�=Rq�`.X7�RB�}O9L��~A85�M5�n�+� *1������@Rh�?%�-q4k�=fӭ������eX�S
Km��Ϟ�$�*��m(ݩj�Ρ]�����$/�d2���x���!�7���=��ڜ8��L���b��)և�ձ��SUJ!�����A�.+_6(�`�_�����w��&��>��?9���2�l�#A���&jz'��>���1^ߤҵcL5�}-wOf�еY�ZhQ&E�aiYx�X`���G�&!�,O)vӈ�'����ƇV���V��i�6��k�T;�!��z����_�D],Y��\11�S��6R]ccr�������A�DL�S��+}ƾq��Ј,)So���'�P�b��`�����"Z�$q����URe1���oB9�����C�o�c�6��\_�p������'<�׮�����!Ш�t���/IS]��rV�d��rڎ�e�pИ��#H��h�Ps��Ov&:�o�'�4�W'�7/�W���3bEh�gO,��x��c{B����!*�lO6��1���x���Y~9���]E�@]��\G�ç�W<�+�㮢p��&�Zk��u�ilpF��Hr��	q�r�������čZ�3䨫0C%����7Jؕ#���n�O��&�ڨ��7����l�윐�S�e�����^�'YI��^=�&����2ޖIh��q��M�>=����Ҥ{P��-�=�Иl��H��`u�t=�W�E�Σ�d]�3HӰၻ���>kgQ�:����`0�l��"�WU�����!�X��H��Lvi������ �mH�<�ú�vk��o�mM�[�G8o��^�̑�}a�Գ�x�p�h�&�nBSڙED��c��:%�.JJ�՗�0��2�8�:�t}�����{4��b�7���=�I@I��87�{"�D��")v��Ol��/�
�`cʬX
PT뤦�H1V���B�����oV�=�er��[WV����zφ1������:@��X�;j����� ���/N���I�1`5�����#?��s�x�73�E��љ쯰{�z��h
�v��.���J���wm�l�A�[h�c;��z��_�>Ss\��Doq��L�v�<?!{G/�Q��3�`��	�B����y��0����:�� �t�\�4 ��6�V��Wn�-����h�ϨRk���ci�IO�^����,c��i���E� ^yX��&��a�çv,�'d���,㸺�">�/u��3���Qp��l:!����L�)x�8ml�4��NAC�F������^�j�e�ӛ%���.m�7���-��}���f����"��Xw�h�;]�r��`��A#`��䫝_��f�z\6H���;�_E^+���҉��h��KzNZ!��e冝��p��?T��kc�hȌ�y�|{øü�aG3�5_	8����Qۀ��[� |9�����)؟Y�
�Wn|���+�����̢5��n�]�%��NHjqӐ��ۄ�}E��%G!�Kk��ܡa��,pԦ���?()�T�l���q���D����R&h2�8n��1}��'��L�}4ݻ�9��k�÷0Zw�z2%�y����/�*��`|t@=��Ee@+)��t*l�F]s���X��� �H�?���+��Wȡ�XP�=7���{�ꦣ�u
�Q�Ċ�={{��� �ɦ�໡�/��c���~��bĐ��5p������/���x
D�&n�l����#��n\{�Q�0Ge�5��b��y�f��`&�3�-S���K�j�
"�>د��Ooȕ��Dy��8��-"�CYa�"߸��������u,�Դ��l�+��Q���2�
wn+PPd��C�����]�Ѓ���xn��q�C��W���_x�[����M�g���]��v��J�-��c��g�|��TI�iA5�B�.e�k�	�T4=�.OPx@����U���w׆ک�r���W��)NU���G��+`���;,����'C����"Q��+-1�8}L$^��<�^��g��m���Y��G�%�@S�^��U�Q�ͪ`��!��6�4�����Yq�Յz`����왎Qs�S��j�q91W��-O��6zU|=V�EL���=ei4f��Ur��p��f���J�}�}��~!�R������y���a{ڠXg��0��K��ׂ��p�����ߧ�u�G�>��_���9�:�-0_������
0������pq,c��#]KL#`ͪ���T.=�G�v����W�jn�=� �+����G�3$���Y�h{��9c��ۈ��r�Mi��Y���cz_�i��g��:|�V�B!�Q�Z�hu6�r��Lᱧ����6{}p�Af�D���4Ps�Fm��%ݪ�V洓6��$�}.#	Pc1L?���@Y�����������ǝ����Ow���GEQ!k*9^#� {�mDn=�w���!²��6�a�#��3�6��.=MV����o��X$kN熅%��ėc-jm��)�+g?�H����-����`�����b�������`
��W'+]�gZ{X#s�ݣHg����7K7���h!?q��!?-��,6˖�%��iZE�&bi�#mm������>��[w����])���_�Si��$����h���&eK?y�(���gm����ӲI�l��m?��x����	{#�)��gMr7�.���g��������� ��lP_䯺� '%�g�&��^��k��N}�u:'y8o<()�����p�XlxVHYEB    fa00    1360��9`*�����f��g�#_)�%iT��L+�T�V�E��y�����!K�-$_�wy}iȂxk�D��{�)O�a�6��K����,�n�:ǰ_Ř��u�iu	�|ó�
�8�r��5��ƨM�k^���0�����v����"댌��v�Vh��цl�9����<=�#��ȴL0�xU9+W~�Tpz�
3�c=��˴�������0S.o�r<8�	䫼߷� �@Nk�В���5� aťC��8���0t���a���2��B��ܞ�R�(�v�٫�=}�@�JI�U4mZCKYJqB����&�i���W�6�O�éZ&ޔNU4��uJUn8���S]-� �Q�����Iύ�52��Q��	�T�M���>NK{��#%>tӔNË����S�osdy�i��_H���-�i/�<����z���e����t�,�z���_FTy�{:�]7f��S���<�}o��������`v�[�e�-����l���!I��;CQ��r
Z�h��D����lx�h�}�A��<x�o�)G��FF��|<ș+5KԄ��I.~]�[���0E7��]��x�C]���]W̩*8-5p�(T���4����Ъ�&8+y�Fb^�%F�#��F����~b<�|���7<&���6��>�%u�05�ym	�����Ŋн�;'�D(���D�	-+����O�߿��6���to�N-U�� :�|��������e���G	��um����p�H�����P��-�9dy�?ĺ�ب�=�7��!n�I�aן��]����ƴ�Z&�0t��.�����wk��ű�3!���o����٤�>����A��a�/F@�4��+5��(�vb��Έ�v �$8�/$�M���᭲IW}��W�w���8�5؞pHZ��$�В�B�TRP�"�n����?��.�Z�>0Or�䀽�z(S�j� �Q?G'n����8�ͯzhH.��Ntt�\�����x��˳��u�b�C<�ow������Y'9U�\�7(���Ag���g]�y��]�G+B0PeP�T	�y��k���P��L���L|�~a���u%�.Oq �/!��p!���"H�� 6H/2���Mu�΂����s������tRp�@Ͱ��&8�<�?����"����zYdBǏ��k�0#'#�P�Z�z�8�G�1,|i(�+2�kH� ���jV�.�G?y 2��8�F��S��.�t���tv�UԼN(���U�΢�"����Z���^Jk�{t*���!�L `�w�����a�x&__���1y=�k�(@Ed�:�;�s!B�|c.��C|T��NM��bt�`s�{0CK��b��ң'i�o���d�r����F�s|WriX�y�z��|>�SC/�B��z4Sy�y��\��I#�e��7g��R9~Gl��1HQ��y3�Q�e�3;Wm�maV���mm�*�ꄲ�Nz.�jB��1!rB
*qJ:�e��f�4�WPF�Alb�;��T��b��u��GF/]5;V�"!GMß��zO�gM�ٗ$�麘���Q�����&�J���Sۂ�C�x_��X��46�]D5����q}�{���
�M9��9��\�8�w��5�s�ԎE�3�7L�g�'��̌G~Ri�h~B�R���7�m@r�&�fEgL7��( ߤ̯l�B@t<R9>̍r���t����O_�o�l�r���Ǎ�C��D!kZV6�Y��ǆ�.�D�)q�\%������Sǲ�}��\c��,�8pY=�+)�T�?����䦇oZ@ܳ�^��v�󜛧�f��ќK�#6�Y��cnZ\UTu�� ���!F�Qy��� �fF���>�wX�_�~��o�$��y�A�P�G<~��~IL��6���}�i$��G�H(�2���u�?���y}!�IUQ��
c�K��p9�c�/>���	�� ��i���Ǣ�Q��}՚#��!����XI��AL�'�����m�94H��s�#��|��>I)�T@K��jY��}6g��݌#�9;}9���u����#�l0@cY��s�\�c��m��ۥ�y�}�ar��f5��6��A��8��ۃ����q�_l�+⑄�AT-Bt}�����΍}zf�d0���!ݝ�x�[�� ;^�)�V^���@"���M�5���@v��ޔ1��#�K-X�,V�iSUq�a�(�H�儘��NC�/`S	3� Q;�a�<���T�;�'=��&�͖_ȷ���F腲ma}��-Ew!񴵙�9��r�gq�q(�!^�]гI��(�--~e�����yk��P*���iʌ�@&�~="[��|EǄU�`�D��s܍�Bev$�sG�~�r����'*���?|g�#�n�-���qJ���X�.�#J4�s���ٴ�1&��S�얝9���[V���Th��ɅC�N����] ��R�n�ݎ��ic���)˪ė2֦�]iK�M��9��;�;������;5�1�L�DbgM.��HZ:[����R�x�8�e���g�c�	��{6*>�V�r�xɴع�M�x�a�К(F#e��Ε���`��>���iv|�L�?��z�:-b'���=��?Jl�,��+H3��/��@`F
6hd�
�+ρ(	�F�b����a�'U�~�&�%��Jh��gJ��; m�f��c�ӌ	{����&�u M-AӺK.�pX*_?�85����&���J�<��\Կ$�zþo8j�y�9]^��M�<-�˃�s�ˈ
�'FG��Mj[/��.
ӵn�m�y7����LI�-�-����\��ddJ$�J ����ܺ��h�
|����ا������͖D bJ�ǽ����e�ᅔ��/2�^�x�-Z��x�5Z#�G-�����q�6���o���>� �I���Y��S���2aq_����Y�����8 ���.=�8�Z)o���o����G^Oa���~sF����e��cE��|�uy,��]X׳���������Hkv�N�ٖ�����@A�_��t�jA�4 �
�:����m�EY�b���^�T��v�DIN)�c�������}�B��u��E܋���[�'��;� ����ZT�v��Ż��?l�p6�A�|`���.ͥ̈��K�����n��\�|01���\yc����	�h�S~�^$���2�r��Q�r�_+�!
�����ͳ?s�"����"��dQ؄�AZ5�K]jn��ZM���Uz7�JSd��}��6â~�)��+����:Co��`b/����c�*�ǹ�0��b�+:]@��q�38̯�F��u�^Q�a��S�[�b����!7zռP�Q�}��@���d��C�M��)��`S�5�XN��t�y��\�n`�} �'��p��V8C�P�/>q��G�"�\�Ќ����j��[:��0ne��'�������.sր��VE����8K��~��K��w���>�a���o�A髛�M���	�T\>��Ly:�wtmo�c�Q|����g�t���5P��=g��^�lrb`���k���D�>����Kf��%~���vٛG-��b&$�	n� .�*�L��/q�<�[UY�T��}褟ћ%M�5�K����3�c�+�>l|n�E�������
ˑ����|�=w
�(mq- �F��	y�l��H�)��7����m�]�٠@@�/:F�O�3ȍ.�M�.�w���'�պ�
��ӈ"J/1.2C�<g�4C�C������_�8P  )�Ȏr�G൵��iqϲX�{_�7��&��F?!l���g�>�^=�=h<�iJ��$��������&��^T�Z*�`����
�9�Bt��1���u�TL���R՛$ޤ��5G#��V��&�1��8�oX)���BMfb&���y��,q����C��3��伵�gRP`������+yY@66���8��^!����_)Rn^�E�XM����1��V��'�7s�IN�+,��C�y�-�j/�Wۂu�����NrU�޼br��.^_�3�Oaz#w�tX-�^�8����i�s�[�V��^Y��v��������28�W&����Ȕ�b���Sʜ��m��L�Y��2iF;�V^9�!<w	O�i�Β�?����8�i��f�	��k�ɝ����q�������Re�-�܃"�7��d����h��Ddm?����� �G�ʐ[�B�_$ln�{��
+N�LB�w�>}W�'9)͓���H5�T�o��U���)"U5ү���	eɐ^v�^��������z��#�>�R>��+Y�A�S1A�6O���|������@pU�W�����(JͶ�A�Sn��l���)���T�I��G]|ރی{*���#~y?AB��%��'���ϣ�����Psw!�F�a��!��\�|�v����Pj
V��}U`���
�����U��M5:dJ!��wX�Y4SS��vu�2�ԫ��l>���a?)�mz��Yo�7]m�W�,��݃���8��{��+���{����u��/�?E�Α,�,<��f(X��5�7��T������TU�	m�_�{_�bӈ;���;
�q�yf� 4=�F�\��-ߛ�!�1�7���@����W�Ȍ� �����-��Pʑ��'ɡ��ޖ6�V̛�c��Ab�� *�'<�P��r첳.����J����wd���A�fz�u���H��o}�mx%
Lq�g8�K�MC)I����������l�ƳN�%��ڇ6�6p{L>��A
������(,j��	U��_!F�Tq-BF�=ʝ�;��-Ż�X�X�Cł`	��7�&�ܝn
om�i�%f�~�T�ks�6��:T����U<�@��Qg�V@�`�s��XlxVHYEB    fa00    17c06s�����Y������.���H/�}����bNFS!�a.J��s�6���,�¡I2�֯/L���K���cF�cvȎ?�.cR#y�
���+&���j�"}N�6�ù��=�n��Ġ��ZV&��c1,�?��(�&#I�8��Se��<5�7=�k���)񠺍����n��CPS�W~�=ĈE�g��^; �p�!��O8Tb{{&G��(ğ�oH�h��q
�.�<$-�oQ���@Nns��a'�V)�I��E�5=�D6�XU~�G�$�(��c�H�0��3=����x�ۣD��մg	L��k�Pf���i���wH,�������^B����p�eHJ��L��G�d݉�����y�}����������Ft5�j_���E��^R1��X�q��M�� ��d������c�%�CP�>�xr\� #P�Nj���(�w�?����mk�1��?~ai�n�"$t_���~fc-�p��au�����6���&L3H��(�M�MR2���,�R|m��L.^x��
�%�/�0�\�g,N�Ek4�S�pW���\��`���-�<��G�+�!��BX�Oc�*�<��4�/��{[�$�]j�&�J�~"�A�[PB�E�)����[�|�e��(���H�
m� 4=��8�"�U���%���oEc�,�k���+��2Ko�o�mW��=�n���M�J�|G�+]>�@5^��K���F���T�$o�(k�ej���k]�K]��<xљ��J�z]�A� vh���7�җ�g6}��`��ka�cl�ն3=��� iQU����~
�pp��O5�ɋ%�vi���ҏg�D�'�17�:��X��ʼ#�~�Ms�����ϑ���%'lX"?\k"yֆ�x�N�_�[�w���ܝ�[�	���}\&�ζ�"�pZw�t��&�a����n���V�`)��.���Q�_SY��d��tZ#��P�wb
M�Br�Z���G�D�xgB]67��[��Q��>����K�����G�+�p�����d'`����y)�QJ9f�?�����(��:o��g�2]�!K�Ie�k>��f�5���O8|rص��0�_���7<˔�w���ˣ9.s /��+�c�f;GB �鸊��:H�D�|laSs@Ē �9{�M=i5��_� e��O��Z! "�}�T��z �.D��Z�b(�M���m�g�9q������r&�_y�	����f�	cg�_��2�X�N_�B��p����n���תh���>k��+eZ�:��,���a�G��fE>��M��w����F��q{�0a'E�4��'*|w'�Jn�y���v�Y���) �;P5�!�����poZݷ\��!�B�|�QzuE�|	��q��%Yҹ�M�=���n�	�.��"(p]���d[��H�ע�nAT��H�1V��������@�ix�����b�
t (ѰQ�  8ը�j�� �&P�I�M�Dزh!���2>*��*������'����ס%��r�i�4�L�+�l\�$�ǻ�+7|�B�?X�;\t^b�HX����B��Ԝ�� -�
1D��0�e�3���5^WX!�-Nzۖ~�R�M��{4�H�e;�S����P�#]S��+��QA�uy^Q��N�7�|q�W�~Ep	�@8�ӽ�~��W!sJ�-t��g	�O�=�"���3����Y���n�׬DY�+*86�$�Ιe�ؔ?C^&��p_��!W��υ.�*��Q�U��	7�)��!�o���*�Z�N::>�f
b�{nb7�0�@�ݪ�
Z�hX��!x��.��Au&�H9��M�|�5��^�$+w�v��~v�q�8!�a���
K%O̮���_�uF2;o��m��aB"�S�tbZ1��+���*�Ҵ�0��/3����;q�4�p��b��H�3��6E����9���4G}�(�^m��G|V��FbT���;)7�k+����ZN�q�M��Y_��q᲼�Ň�-smPnHg�ː�O�7'i��K2�O�R���^�
p؈c�A��O �uS�,*��۱=[�Z�
��{��]��E�͈���IV��KT �F=,�z8����^L<7�cݵeE�M1?�	�
t(���>"ӥ8=D1욎�1K9�d<��� #j0�6�' �__I�!(醦���'�������a��Zm�O�EPbg4�^����)�jB_oA��Lg���*	Z��T��epU��LL�k���"���L����{8���0_'(���j\)�+��f~����$fQe���?�>"۴@cwa\�.�h�̗�oν��qR�'w�zJ+�T�7�6��zJ�q��i�K�E�lt�IXB��w��3W��#�'� ���{�+S;�q0n9vg��נ?�5�9,�����$�P���Y�gvw�hg�b��.2����%���c���-�}7�ڣ��\'�W���L�G���s��� ���%�:_� ���L"���3��Ar��A#��	����5�A$��S}���
\��4|�)�F�s�\����4:�3���x'�t;_�L�R�$[/��*��'L��R��m8�)ES[��9�g��ַ|���y*`����2��(72�}ס^Vke�3�hF�V#�m�c�:�*�^Җ/\�I����Wma�*���,E�P��ev6���j�cX�v�Z���6�ܴ�N�;p�s����@�k�:�g�!7ޏ�E|�����n��Uk�t�����a�F��3d��pw��w6Y�'������o`�d�b��z���[�B��oc�L�[���V7�b��L��\�zoԦ>�PZ6���C
��-�b+�o��������J�K �O��T�;��+�qZۚ$%h��0ٝ���ǿ'����Xm��舋I!�nD�_�:9�X��@�,a���y�����yP�ܧa��u:g|pp�Q��~A��D��P�9(C�I2�n�y��h��*��<�0���!V�>`ŷz����h�3���|��2A�Y|�O6�I��Y�'`Ya���Tv�,��"�a�e���ȑT<N{�F��s}ɪ.��2ws�!߫�)��M�q�$��l;�Y��(����$	�AR�Y�;��ł'�O?O����D�@Ơ�:�����3�J�7z9�s<ܒP�\ ��-M*bv!�t�/�	��_�G�ʀ�̀ vBOe!ظ�ޠ\hx����~K30��rx�x]�϶� 9�3iWM�yOB@Ο9N�����Ip��z�����e�ɋ3�L����1���c��A�ۑ7������ܰ�P����N3nu [6� ��qR��&���<p50��<�����de9��PM�O?��)�a���c�A|�"}W�Ӹ�)	���*���a���Y���0���}ҳ=�`7H��y�,��Fx�g�̢C��ZV�>1�(K���9�,�ØxZ�Zo\�wO���b�cx�j�q�gAA��ؐ�yAgbk����c#C
�c���I���=v" �fl���̓ۇ���UcQ։��=V&�ձ���Õ����l�M-�ķ�[^"�8=���KVwg��
�}*�#Q��P�H�����B��i���ګ��'�t�xH4�BV�P%]�L��a���7���"��[@���"��^�8JmE�;�� �K���3�g�=�E�z���8��>;I[�, Y`�����{F~��l+3��O�u�y6_�l�6��s�������R�5�D��ۡ�IN�)6NH�2�L�C�����U\��V�Zw��I���/i���Զ {{��k���8��.�ĮL�Q�z~-b�"���Ly�Mb��*<�7��_�	��xm]ѕ:hK9h!�����e=�[2J��E _J���:�עە�gdE�e�p�p�0��P�[(�&����bld1W������D"]M�:���M�5�b��k~iq��ݭo!���l��2
�"}��?�9��b��z��
?o{+ݙ<��0P���N�8�?+O��ء��E���ߢw�awkCc���\�3SӰpb[�Q�_��j�n�dBZ-��|j��L���A_@�f���U�7�oW���-:F������v�S����Hb}G�XZ�f�Gfޑ�ü}ϒ���v�ܲ%���R��W�z$�{���=k����VӳTF�~�ʫ��<�O����ʑ�t�v����Y�y�������NA�0�2�:Gr����w���)�����q���_֡'C�H27�Z���u=[�Z�@���LY���y^��1!�w�S1�-��E���︑Nʄ΍��EqmJ9��\[Իs%OWi��)WĶے d�\�H�IvE�^�V���R+��L+M������o����W��mj��t��CR8�����\D��m�� �s��;���]��3jN�N�$����<xY��� ��Z���<���� �����%��&P��A1"sFb�
l�.(;��[�dM�7�$�.	�ć����K~Wx��#m$N��I�{�'�/�M�7�{$��c���$������$fi�X���F�	�HdeOCK�d�HZ.bp��5�ٗ	vHtr�柜B�A%�
��,�����b���Q���b�H��n����؝3���\�,�9�aW�z�F���d�fa��u0��0����2��zl�����م�7'���a�E�vWǞ>q���'@���K��5����=6?�t>����r��kJ>o�g�	�<� ��fVH��{ώ-!��Ә�:����P=���و�c���BK��p�
� ��mu����6.���A�V�K&�S������beCr��q>
M��c�GG�?�Ƴф`"�Ƥ�~�w�`�׶�o��ʢ��7fS��U��c�D?��V��Rv�(�i^�KZ���0,����]d�N��S=1�d�T.�������݌��QH�b[��x?y_�dRD4ˌ"&�6�yh����𨪄����tX�ѓ��N��ial��,�I'�	
�s[��t��LO@��^h�t�3����H�L�A�4Җꗡ�Z#Z��N����*@L-`�=x4���9���6|1t�����8���oVu�G;Q<g��%�P�6��p�-)Z����G��U�k�6F�X�T	7|�����L]��n�q�NX<����L�IҜ5��j屌Lt��-�$�w������e�GY������9��r�㱛��c^��1��� r�T�X�/՚����L7%�3�Ka%��3/r��b�8�(����l<��9�_%�`�4Y%�G��ء��i��(Vԩ����I(4������-B���8�Y���ӳ#ܻ޹�Ԯ�Τ���]���n:����'Z�'"0���Z;]ş�����2'6�?��*�J��p�'��i�i��0(��t����Я�&�pw�x��e���Q�L����V�c�a�S�P�88-�w��F�Q)��n}�i���ߎx�A.xk �6X��f��r�ZSX�l"��Z$K}���"�QZ�{����%��H��л�����l>5��Zk��1�$�gFI��<B;{�	G��d���'�&����NZ�w#��;���-��})2�:���qƻ��Ѽ�@��ӳ.rılKJ>9�>����ꋖ�~U��9"��!f��<����_�/�s��s
�!��k\������rZ�ϓ3��]
!��?���?!r�$&H��1�2�e�ş��X}��Q��<�:%!ޥ��+͠�\�:�ij�8�8�d=�@DR
�is�����6흗$ep���Av��L[Ad�&�1 4���u>0@5�[R��Ȑ�,�c����	+�+ b�'z��%vR�:m�%3��b���:��fa޴��������\Ð���-$ ��`�_�s�?�2t��W�߫>�U��2x��(RW��v\����eԴ�!0Q�W��p8XlxVHYEB    fa00    2290��t>n�m������scX_��dЃZ-����O�U�v*�3�=v��LT�\�� $c���uf�EHHҳk�kJ$��~�Q����m�׷XĐ�:+g�('������"ۨ^��;�
��� �L������~���x���+?��\����Z'������!�C
�E�874�X�����r��嵨P��`��p�Lt��ڮ��{�&�%7�!�h�#���Ϻt���=c��^˞S��Y-(�-M�p��6$��@]�����c���D�If*�� 0��<p�+��׌xD�'6}U�1���,�`J1S���I�B��,�Bp��9�����[��k��m!�QP��3G�kǥe1�ܺM�N���R��×դ�Q�|�Q�LC���bRMï�~�z���5d5ꅳ�RB��$S�8�����`��|��1�� �72Q
���ܱlڄ��Q�2�9I��4F��=-���/0��Ҥ2�N�&��|4��c㭪���1�e&��Kɹ��J��UcvC-���͗�_ZZ��/���3��.1������k����H����8I�M�2�~`�;����~܁�Af�����IwT�3�@?Vs�����+���{^��ŷ���uIP6\pn��0�s8�Jم��#1tz2,5�.6��ێ$�W�n����؁�>��ւ�P�r8�u��|݋h/���b�5,V�����	j�Z^����v���|{rHFx���(�UW[�JE#���Ћ9��7,ᴙ�S�{��%�Q�v�Z_���A���aS����O�K�O�P>��[,��$��W���m5XHC�.>:��;�D>��]����PC����W�.���m�uK���J5-�UsN��
Ǹks;"�ܤǱu��Ҋ����Q�����ް`p��j�B,kku�qA�E�^��;�t��Q�&FE��T�~���;�z��e`t���m��h\�h �=�'^f����/Y	:
�N��ʟ��W�`P]@�鎴/6J��?�����\�F�:~����'
pņ �d[�Tڸ����r�y}�S)&Ɇ�l���������'�N��������C���6S$�Qx��ε;t)	;n���8�W�պ~���6`�����GB��4R���aݞ�'=��B�{"NB,UV��� ��#ψ��#�'� �h?<�s`=������]��o��a��,����\aqVY�W}�������O�E]���, 0�9��p��ț��E�%q��������v#)�M��u��4�pW#3+HNH�0�vm�;�o�l�S"�R��]�o�c�/��e��DŮ_����������7d^(��1�˜��~��Gd�tP�s>��<�e'}��nU5����3Tc��[�e���i�t��i�ɝ-+q�Um�3�,9.��Ø�X��C�w��(i���;B|j�b���̧�![��m7Ok';��^Q�;Z�"Gf���JWp�eP��.=�B.~�/���YА�����*rW�3G��?H�����ԮG+�[��4�(�b����-3���O��'�W��ay' {F��h��J�kDl}p���7p�����o�f��/�UzK�ʁHElǔ�O�dQ���U�D�(�l�Zk���z��޳�@ݯ�j�I�<$��	V�}~i,����FN����T��@���C��ok��y���f�z��H��1W�wy|jN)#�X����؅"P�&���?@���pf�_G���:߮UD���*�:�5�	s���	�Z,� KE�4#G���"��H$`�.�ˎbP����̔11��4���hS���^���$Zl��p��4�3-�>�±ؖx؊4��s�B �>����������g�Nz;'�:��N����9��a(ǉ�<.x����[4b�@b,�����W�sJ� K �+X�1�U��Z �L���;����aP���!b[E4vtQÛ�wP�����K�c h���C:cU�t)5�h�;1�\����,<���6�N�k^��"�l���yu�E
�N/���L�G[��n��H�����b���&���^m,��
��ɻ��ɩ�nU�-?���F�A�N6h6�!��X3���~���F���e�+���DY�*�%����BHKJ�U+�� ��/�ZP�=��hf]3�D)�2!î�����eW�U�w���e�v��(#�.`�(0�u`�ͶG����L�WWC��G�������췭{t�9~���w����r�]���A�A�&7�>�=}U��d��F��D�a���ɗ��P�8�/2�~�:[��$�4)��j��($��$��=�	Ja^J���iL6�<�:]��)��j2���M�L�$�;[�V>N`F���Is��cKd�T�g�{�Mȁ��lH+%��M }�D��؏�*����)�c;�'�I҇�:���ǒ�(�M��w^��:Au.#̪����$�$(���|S>���\Y�P�����ҤT��5Q�=���}g��8Y����z���t�c�˯@)�>���V�h�1\����C� K�z��GO�(��1���U�4B!͜=��!��^��9z�0��<���N��������;_�����;�2�������hn`�<�-����r��6>����A����MAqJ�3��ڻ��J�
����/����%EY�H�_g��,�ֳ���c��u�/�c�Y]�#?�u	8 ^>���k�Ax���)�gOy�hh����b��'0�駈���Ɔ��Ɉ���Lɮ�辍Y��87I�AB����dm�:���������!_���d"�z��Ò�&ѬU�y��C���B]�����;zn��W��G�C�ш��@�ք�������%.�u|�tf� ��j�_�D��_��z55�~0"��+ly\��f[�a��U�(�3��c���P\� ����-��S�K�(XYVs�X��ך?���9�W������=�ߍV~�]��%��U�l�����#�����:I�E��[�3MܤB�Ba`���f����	�����67_A�i:����ǵ��|2� �Y�qa>�[�,8��9%�E�rPp� g -�����0fz]aT���s��a2�q�ʜ��	�S5o�\_!�$!���
�!���`|>�C�J`
��'&3e��;�l�5��7�EA?a�e��k~0ӪB-ʽ��a������6"y�M�N*�"ӚkE2Da[t�;�۷���G���Zw�� �=a"_� �6��ߚ����=�0���$���~%B32��oH�p}p�/ֶƨ�1����O�o@���؃��LU/�q��^�8j��S�����S�X�	1�\�̨"�C�@���jp_7GV:ˑu��� �o$�*��F+7��tuR�"gX�_�x�zGO�� �)jd��I���]}CO$r�{��B�m��ox�D�~*���uiNv��x!��6�[P|�Q�-�My�z6Ԧ��J]9�Dճ�@3�3�فJ,��p�xo
a�-	�"
�X;ՙk�m\��#�'`�V����}l��$h�u�S��
��%�Ϳ�!�[;���lߜrl#�'��>�A�H?�Ԑ�k�;�P'�+Wl��#�1����{�{϶R�j�`��Tf�2R�2f���i+�x�������Q��c�luժY�v��6 ��;5.X(��L�{t�f�h�0�+o9�Le�ݻO���ˇB�-�b�����{����U*�+8����m�HI ���%H`�`���˫����b*ɨ
�!�Ņ��˧�5�z����y2��3%D����M����&g����p��;���s͖	�B�M.
���$X6�ʬ�Y�����<]��a/O^��.��M������G4�*����y�IXl˺}�ޥ�HBW�*7�Xk�[��V�g}��.U��5]M���]��H��s�m� Qܰa(�V��̞E��>V������c��Hz���M���i6hv�w��|^e�V���)��琜��2��3�L93��&px�*�b:���Ώ]0Xi���Ϥ@� �ٛ]ƹ1oP>��=\��,k��.a���y*R���c�3[#�Vlgv/���+7�{l<���!����΁��C]�[0Af:O�]�q��)�)���ߟ����m��ByvLh� ����V�̸� ���<�.A��q�?ه��}�m.=�(�G�L���~}��@�U�%��U��=2˴C�6;e*4�yȚ9����X��rJ&����R���N�K��p}g/�����U!��<�ǡ�dTaz]NK���+ɲfH���k��9 �g��ͩ�Α��n]9���A��&�oAi/�>c�OOFg*����dY���ҙ�AI��e�1�D�����fD �fI���X5F9蟉���Ҳ�$Kz�f�٥=����t5�0K��g��&��顨�_$Ǽ�� �)�nĘfx#f�;m���rkҹU��C� ق�G��w��+,X~����-��>A�F��>[v����D������qI�L}+���X���8�۶<U2�2��9P~�X�o"{L±`C>,�������%��D61!sB������yDP!��z"���K�U�\O�ɜj��gif����V6�8
E���Ȱ "(�@�.4M��;�%Z�y���X���}��q�l�A���1Pf�k�Q���5����d>�뎌t���z�>����Ϲ����=O	.��oCǎ�ٯo~C0��kg3�P���\q��Vl�Km�e�4Aq)��� ������ �{\�>�Sg�σ�3�[1{T�S����qa|�5�	 �{V�W
�Oљ�rh���,K�(Th��,�������oOis��#��n��uq04�� �X��ONޱ�R���b�@~ԕ$Bt� �R�|�,�g�~��6��ZG-:/�9��7�
џ�8R�-y)����Bd>�En��,}���� �1
�C`� ���{ʣSk=��4@�FK/���dMz�߼�X��_Z�!���4<��C��g��u�=~�#����af2Qi���%��ث��µ�wl�kIz*D�#��z�Z���,���U�͊(*'r����ܳ��@ya��|{At�0뉸�nhJ�m�Y'�� ~��r� \ek�j�f�*Y"���*�����n�!}F˧��C���\Xǔ�2M��_�\��3o�i5�a8V;"�2�=ll��l�P�_T�`�G����:��m���Fд�騲�v�����w?��偱�yJb��m�,�J���Y���?��$�ofp�S<	e��˯�Z���C�8���v�G�M�ݷ���F/������i��i�!�n��B���C��W�r�(dc��8b�&�K1��<�N�7T圐� ~Ȉ�r����$�/���ҊSZ /��3�+�ł��j������ۣ�&e��\"\R�×��ܯkx�ҙ�~�K��&|K*�I^R���c�J�#�Y�8;৉
�E�u���Azj$�C�`-��o�h[����ih������5�E�ۣ���s�@񙬩�u~��jB��j]K��k�2mJG׿]���= �ؓ���0�5�<m\z�?�ou��pX̡'49�:n�#����Zh#�ڲ�	��?�����3��֕1�5f�K{}g����@�t����z���8�kP�L�N�����J<R��%�k��lT�k�x@,���ć^(�2L�AC��I�g�r��7�[M`�#ƥ{��?kg�7��ź3`#��R]%m�����|�Ǡ�.)_��&�/�'��g:������0��l�n�m��~�{hq7QgpŃn{V���F�G[�7N�cܗ*�MH{`��m��H}m��)�ǧ�x�ڠh����{Z�@�,�%#�D����ݣ�!�^�ySok�c�3M�����v�L,G�t�pU�k�%�#��1� K4g9�*U�I�Q��y�$z���<,�_�KҼ����H!8�t�xX�/���P �>��K��k�E6M[�ü��ِ����w�Y-՜5��f�~�f���{�zO���6 Ƞ�I��	���4�$D�{K��s����ǮΆxv� -8�Eap�5s)���.�נ�#	�����16p���)��nCa�[a��l �/LT�7��i����x�ė ��c�-�d<�@��Ù7��e�BI�\��jq��#	��:�C~�@�x���Kw�̔�S�]�53�)9����5cM��5�Ft\�[�<� ��X���z�~�a{�� �"Q���T�2��k{����a�@��1�����&xڄ�3��Hn�	��#֟vR��[�'���'T�J�F��@�PN'�w�zH�)�Z���F�b����8��Ʈ�����poIn����Zz�/�Lk���[I����N2���XG���@��k*[�ƍ��I�U�Ó%�da?�V��b�D,F��qs��X�5 �_�;�Zo�8����釮5����̐I�Vb�n`C	Z����f����^�03�O(~$�9��{���$�V�0���7w�M	������S�R/��X!�ؖ��m^+T����s�R�`~�J(Vtz�z0�*�9�16h/]�'��.�g1�`�8$�����u򩀔~������1�/,���Ѻ�(:an��AjE���)��m�H�j�X�g<�Z�%P���h8�C��_���6�O�\?���"�0<�'}�Z���/	"��(`1��z��Wv-^��FY�ga��|\p����W#�eWR"�3V}H�E�+��\�����)� X�G̀ )R6M�u^0�{6��	H��{��G�gǩE���j�V��$iL���^.8��%� ��tN����c�\3�vS� ���iq����9Xw��!z}��am^uN/�~(�zqi}WgLo[��8��7�]L)q�p55�AL4r�Z���_,�m�լ��J�&]
���l�T�-�Zl��)�ҿJ��J[�易cZ<�g�.�MC�����3tG�k�%��K������n��
h��KW������1��D%�0J�}�R��-\�4��XS@,X�y����k��o���Ny�V聸���+��[���n�TN�3�[s���vve�������#('Ɋ~XafU����֘��8~�=�&j�m�2P.g��/�-o��a/w��LձCY=$����C��^�|FQ�$E�%9�]H]? �o��u�P}e8�x;�d�p�U(�o�ڲ��I��t��-�jS����bז����K�e4T;�����3�& -�s<�5<
"���4a0t�˙E긷��P���ka��̷�(���Ua�o��nś �]+|�aAw�� �oIZ����+��BJ�����*�]�kH(�"�E����)��=W���9
�Σ���n��Yd������o�@8��`PD��F���O ���8��@�2D։�b[	:�`��F�L �IPbHiT;��hz�l!/F���W��7����@��IQ�|͖���5����&(C�
x�{D��L,+�ّ	��4�3g�G�Ap;V�J4����YK�;����/�������in՛���u''fؼ���=�v!\u ��!%��CY )D�N��!�x�w[W(4֠=̰I6n�D��9	=F�'����U�1r���lB��5芿t��~�?I���xw2��o�:��T��[ɍ��n�Vv�"$'k:�*T%?D9b9��>�q0��j/��8Đ;^ܬ����
�8Z�����>��������ϋ�����<�:�$ܴ��d^BD<ZA 1ywx�G~j䇊��]Sk�ޞf�Z}��uC��x@7�E��'�!�B?*hH�穈�U<���v[w�lD�y�n��?�
����rW��ĝ�FoZr�!����)�EuO� ���\k��J�m�/��1� �Yl�2� ���k�z޸����ѡ�E�&;fg�(({S?�+��/���(5 ծ�^@�ފd<�J	�~�R�_l�,��-4bbݜ��J�M��"1�<�#u�WƆ�<����qB�(�'�b�RA�gЭ|-����W��O��NO�Ҭ�*��L@���N	��*�<�G�w���󏫂}�+��Շ�pr���J�� =|zpld6�D����0��*J� s,^9��y�6�%�'���K�-��q��:$eem������<�gi�c㔵�a-�[�+�6���e�2�\N?��wA`>'�0Nel��J&��@����d��k�gR���
N���})os�K���&*�i2.Q�˾�V�Mu����6s�\��'�Er�O˰�<:|k���2��RS��=��C}��ޢ]q��>M Ӑ�=���D9�{��V�iI4�ZAt�^��U>ѹ�t絏H>gN��i�;�[��#�3�mX�L�l��h�M�Dy�����J
Y5�n(!�$�,I|�;�C��(���MŎ�����ɥK�wQo�]!�ĝ��<[0��*SE�շ�������?�A5�L���[��aѱ�ȇ}=Dbq��D��[��.0xͱT�,`	�TsØE�C.�YF�I��w���F�rf�W�ē���q��vD(e��ԬK�� �gI�=����� dEd��K�{N��5�z(%?j��ϝ�{OXlxVHYEB    fa00    1f90�J)�z�_ATd66vZ���,	��0��S�2J��m�:܃�w�( r�U>f�r��c��j�� �5k�c���*Ha_Pľ7��' � sWL�-j����y_�vk!�mq��/݉L�ƀ碪ʶ�i�͓6�W�>C�M�f���-Ͽƻ��`��V�
7��4�&pir�DX������t:���,����*���פr]�+�b�o� ���7L_�f���8[;��B��PK��y��l�E�t�����~XrK%%��­v�^:��W�V2�����t�DY\��� ��,�b�V���߹���\cR�l���m�\xմ�O�=���Ӛ���P���a @v=�pI׫�4`�����])��dP��P�S	�e�/��,H7��e�Ñ���������a�1�.u��`����̝����Z,[� ��FyT�X����6I����tw��*�)�
��O�Y~�j��v���P�����1��2'�������>��ICD��c�`U�j�(�xUl캨�ak
�xMN�(��G�|�B4�#�m��Mlm�Uϙ!�@N?��b���5�j!gC���+��bM�l��\_ ����Þ~@���.�|R���X��z.H,AQ�f�*�ur&h����p��P7�UZ��A�lq��sM�8����R<�"=���	�� �L�h!���y4�l3/%t�Qzo������̖݊d��y��d;'� zd8f1{�$^�t�ikH�-�妩�J�,�?Ys��ڻ�7��G,��Ƅ<s"��W��|>$X���'\���b<s�� /|*�dJ�(ů�5�v��eH�π�<�ߥ	_��$2��!$�W�p1����DH�5Ax?U�;��������F�sIF���1�Ft�;$yN}֧Dq�}dp����B��H�Axj�Z���c�#�P��vgIV�T'�0Ğ����|g��M%�x;Ge�\�'{�%Q9ݦ��S5�sQ��J�^1�l�]���`�\�SS�&�ڹ �H�	O��@���-Ã�R�
����&��+Ҭ/z�ДG�m�n�
�@�X=�-�šZ����kr����m���3d������%J�Iy����\�{D��s�隿�t�����4�C �6�'L�w�=HNԍx����([&�t��%�Ӕ*��'Y��XjJ_'�� ����fN�,�ހ4М�`V�o�=i��,�"�Ѩ?�\�����3�>����M:�`��RLIvr1"�X����ɈI�^L��\{���:f�����a��}jl$����"2��(}74�Y
����$��u ��.�V_��%���������Lo[��ח�Ya��媠�����|��;d������[8��n. wL ��yȝW���Ɛ���C�&�FA��qH�|��$���{$�_�t�[t�m�2x�g.tI��N@��[��������8nP� �j�`*wT�걙��f�mP���~��{>e�ʠ��+�}Դ/~�܈��5��AC`0I6Ye*u��9�f �=���N���Q(X����S���� ڰ�l}f��Q�+� ��ʒ�L����3�5�=��ˤ�B_Zٲ6����Xs��Yc��A �;�Qw�G�rYC����0�T%l�z��i�~0c�*��(���Ά�l����98��ꛐ�n�험�E�%i��ז�k=����dO�%���0'�8���Q-���n�f6�|w��~�Z����*�1�1�5����no+�������e%�K2"â%��n��q���NH�#�Ea
X�{�s���+�Ph�lA뱪2]o�7��2�߄$�2���8��Y�0J�ڂ��q��(H� ��sC��3\��:�h94{�$K�Lŝ�k�A�Q��7F�znֈsjdK(��C<���?���(�xbPb��H�8�� K�o�f�i��td�L�MǨ��bi2w�Љ5:!p]FA
�m.qI��"��뚊?�~����ݼmF91��v��낓w����QUQ�� ��(����TZ�LT����4jY� }Ru������1��e�f�2Y�H3�{d�CF۹@2��f�U�BU|�%a���%�U���&L�����$�w�)RP(Y��?�o����o;�($Q��W�y�Oñ2&�L�(B̰���0:	���<�f�mDl�	�Pl+�XQ��]/������u��c�b�/*�+q�ߙ��4�e l��@�# wBO�i0V�4��78�]�==�b�W��(ezf7�1�ڠ����씬i8.���z�r���p/�n)��IlwI��#�gn����+Y��^L|��<�FP>�S�G(���"i�Ċ�IZ����d��Ϊ� c��E��22�D��"�j" �7 $������-��z�|u����M�o(���Pڳn���8�|$g���9��M�@�c�c��S��cF_T�
��;��K�Xbm�d�3p�M�k���������.�9�&���|m�3���~[�n����V�i���(`��sm��e��7j�*d�_������>��_��(r�L=v8�E�!�:��X��jo�W�ГU��k�+�-��1m����O���FI���W²���8�)����s5���7��W�#���x�zgk���_3CD�"x�g���V��T)X*Z�[�O�����y0[����-� ,-d��H�P��£|��f��/��8u&R������v�l��t;H�X\v����h�zQN�M�j��D����D/!QO�͎�Z�.�<�~f{$���]�鈆�t��e������>7��|z��p�D?��C��xW��K��9K�+�J��tH�����JDS��GS.[s{k����Ђ���O��:߿e���������\d��Q�����W)�BXl�-B�%��*�=Pi�KRs�R~���X�p��i��8U���ii�	�o�Ĭ���H���(P�����{8��K�]w*�Y� �<���iK@N��أ��ƥRbP#.��6��A�2]��w�6�Eό�V�/~�[�����K�g/h(�7�+��[�$�A��o���L����{)�\J��K�I6���'ִF��K����2O���$�oΫY�xGYKg��JV��5;7$z�q���\�@��y*!���x\�.��4�#�����J��y�Q��E�cZ�BsD��Ap�"�ؑt#}���m/B4¹a-�ugW.h^�%�ȏTZD8Y�����6R5[%�P�*'���$3́Q��w���d�QqH��t��C}O&�D��5P%؁�BF��m�������v�����;��ʀ��E$�8�:9$f�Nu=���
2���9ϘY�/�E'�&�Ww����P�A/:�1��*��� ���Z�~R�6\��/C��ð��8��X�UگD�ď��qB��e_Nj�qfX]���Ő|j*�H���}jޕ���Q+�֤�� �NN&�0p=���y3ث�y�Mw{G��M��urS���į⎜�1]��hA�d�4��A���z ���eU�W,�I޾��Q7���@���qȞ�Y������D�6����=!4��뙞'�c�Fw�3�KL���|�\1��L2.��|�Wm
�e�K�RA�J���^�и�������85��\�Iy��P⮪�����i�K��`��
幍�9o����|@���U�{W��]�Ƀ��G��2���zDFyD�!�x� � ��+�2�&��(k5+r�{CÀ��k���>B���u���j�'��n9P���+7)Ά��EW�uJ"�2i��	��(��W?0����)u,�N��x�&�~� �b ���*��p�mT�\BT�پeG�ś+_v�ɢ=6���q�����b~�\�].s)�V*I�t'�[�(����~�%N��g<;qc��R�^xL�\���Y%���kK��a3K�7�J� �vOŞg gv]�6�bG[��R{��������¥�yk��_4����?��� ��a�Ù���,���Z���ɦ��_���05��]��~��:��**M��M�j�l�{�5��f��L	�a*��;�	����+�|1�X�;i̓��Ѿ�����8-�����c"t���&Լ�F�����8w�2hJut�`V[3``m���:%Y���Io�!�4BD��v���\\e����K���V�� �#ҏ��ż�s0�Ӿ���8��̈́�W�^��eO{Z�:���Y�!��~�)n3�_�^�Y"���^���@�F�-��c"�v|z5����\���_�/��݇��gnD>�g,���3'��p6^���k#�}�7��a{ �BQ�DSe�odC��Ƌ�H��ޯ��R����A�Q�5�(�#ph_*��7кi�(���o��C����.����J$������bfcnR9ƯՇS���z,V�V�ۘDn30�����vLģ-g�đC�s0��?Y��X�*���#�e�8-:��)����>R-vM-��FhU��#���R��)�\m��3i |��랝Y�����T?=r�r��^�ƹ�u��<;�R��2hoz�R�	���˿4�� ڈ?P�M���K��ptma��h�{U*��4}/!I� �!VLl�n���@�l����:�6�`L-�X;��'"}����O��!���l����B5��=tv�.� �]h��F_��6΅��&�h��
z��rAÍ�ûs���ky�C�L����k[�夙��OmT��,i��Ӻ��wR��&	�VZ-z-�E|,���?hǂ']gN~Ѳ�,�;���V�˱�������j��_kv˝gg���ʊh"���^r#b�����q�G�Z��w��5�]qX�n4�L/J�����|�k�<�$���^�׌�
E�7z*3� 'j�y���T����:0qfӱ�:d=����h�jw�ť�I	o�Ezt:1�D�c**��ҺNO[e�����6�*#����A�%GR���mt����D��k��X1vm�R)J'>�L �%��v.M�jL�q��ɜ38P�|&ۤ�gV�i��7ߛ�,R�s�F�.6������{^ �#n�ΠR�on�.��`}��N�|�k�u����3�!��g-��`�j���w��������2�T�j�Q�,���l;�Z}q
�-������{�)�I��tj�P�2�E2K��9Q��s#}��-������&��"k��D�6R��a��n�s۶FУ�Nf�5|�o�ES/����^̽��?���4�x�p�¡P<t摈��nMm�t��8�D�tZY-i�Z��Ht���U��8.p낊�,�4��ս���.�N#B~u��!��1 ϖ	d�����9��e�`>��R�
ƹz9�d�Q[y�/=p蓧���'���-6]���[��T��@hk�U��g��kկ��t`�
�
����pACv��|�dT	���n�'��,��Y�1���~�|�e���t���G]����L�aUCӢƪ�^Y!8,C��W��F�ְ��My����#�<w�9��z�K!��	I9Ő�U+�p��Ì���ſ�X�f�
F�q~{"i���w�%	�'�Iie�5yL�_5\�\�#k}
ɉ4�¸6t{��3�j(R|w��
��р шQ"��=���\Lݩ^8��-�B��Ģ�^�^v��-�a�nom��C�?�<D�Q����reL�,�J6 D�7핌#=�a�	@�L�&l���<�g`��H�9�d��~)҃���6�X��	@4G�ˌ#v<>Qj�H;J����edU�ⅮYg���l ������'���1?��;}�:n!��Z=�TL�~��[�*�����|��-���;����ut�J?�U��T1{NV��h�{�)�M�ӓސ���f")5��d�A��p��6�NkSܿ[t6��AA7��8������<m�u:"N��Z1���bo�O�"���'ٳ4�H��:�h���Ѽ�HĘ��Ҋ8�[cFФ�6�ڤ�f9hv�Łd�ͱ��=��::4���L*��bsH��<���!���0Q�L?Y!p-o�I�,����.w��R�����ڻ�p��P(�.H�����.�gm(�����m� Dɜ]�>�1/=[����x�"�w�T���!（�~����a3������%m�}�	dH��%WN�\���R4�Si��Q��=��PC�wέC_�P۵Sdfn��.}+�j�0?�m��(�ea�P���2��<;���"ظ���H��>���_T���̼�(�6�/�s�c�6I���Kn�*G�$���0n��+F�Ě�ꏙ����;����8��PRLJDT]�ςػ���'(&�½~W3U�,����6��s����X�nt�O�L��	�1���q+E.�l�l�qBC�냆.��֮���Y^nxrL\�T5A���o	�d�j/^t`ӴkJg�h�6l�C$oP*���gZ �/�F�4l:d�e(VYz��hnD���`��_6���Ϻ�X�jA�~�'��[�,*�}�}��D�~����f���>'a�:�A��睲�Y�����fXl�'�aJ-�w"g�q0�Q"`��iɐU�}e!�]4\G�G�ؤ�ڟ�7��\��A�f�J1����u�Z�aP�@pp�O(�J3b��b{�fH,��X�$�.�v�+�+��z��+8��q���{
�V���0�|�7��R�V&�g�i��Hto�:�����&��]�k��W*�5��!]l�9�:S�x^q!��#Q@�'������c|�9�$��/�6bue	�f'p8��x8��=v�F�UB���%U+e�� GB���#4���j�{�4���Y?��o���;�R�x���4���Dz/	S�̗�������B��͟��V��)�ཪ$��Z��O���*��^�a��A�p|��D�"ʉolõ+,�pp8�2i�T�<��	�S�`l�4�`���ۿ�E�~^�'`\+Yq�!�
O��iR~gGT3C��>��~T�{��e^"��r�����U����mõ_[�
��n�zQ+MI0u?4Iq^}�wq�鯉�2OW�Et3k�w,I����_ҍ�vd7w��e�p/
��B�i��Rꦿ��'��z*�	�F���3�X��-�QⳈ*[2�<�_�8=����ӈo��<D�J���Ѡ��u��^8��%��8b**[}��-Q��oY���d��Q�f`F��%06 �C<e�}} �gKƆ�j��Z�+mM@��� �X��b+|�7�]Y��u��σ:�A,����!��`e���\�Ы�HB_n���h��S:ľJa�,��w��_d��e�����A&�np���>!<����Nl��$�ƓӞ�n���𘷚Q��x�)FZr�y	��Y��ݫs�yS����tD�#a\fz,��-�:� �*�;�^�a�eg/�D�RX��>�e�ƥ-5��*�ma$�w;O`��U`޳�S���	֩�����<.��w)��u(���yK*�����--z�,�9�V5 �8�<��
yw9t&�Ger��AC^��i��G����w�;���0,����x�=��Q�s�WQ���Q�e��;%֊u�xJ��'
����-�f��:���|<�=a��0�U �sH¡�8E��Կj391"�ka-D�!.����'�W4/;z�T�s4�����K���}��! f�"����Cg���ٳ$�eh��>6B����e����W�2H�; Lj����$[�h^��+V/�Q*;A�q
��D�@<	��N0�iܔ��T {w5�C�NH�
5��7й��3�`}=�sDU}�#/�h#-<�N|�}Yv���m�&D�3�W�F�������Q�
�?��KvR!e���"v�!�~������8��v~�D3z.wz�#�k;��^s�C�g祵R����aXXlxVHYEB    302a     610�z5����C������q�~��MSg�d���Dk�j��/M�p�-C�:�b(�h��p,o���I8�����U�&���K��=���0�m��D�(�tnӲ��J-�ظ���J���6[���8���L���H�(�]�fm?�X��pm1���%��]x�D�5?�OiJX�!F�t�(�(s�7�4�.C�4�lI�a���9���J
北xoPV8�1O�<sx�q��=�x����9���}�kD$���I� �O�eHI2�M�����
�y�2���O�32~LC�8�=だ�^�˖�怜� �"�~G�<����Cת���GH��f�,�(����~�Wj&�iM�+�21��xɀ�F����1ʹ���P� Ey������a�4��kZ�vr��>5�׻�������ԅ��I���9���Q���4I�!`���n��+� (��N�A�hO�ٗ�`�2p�E���@�p��=[��Ԗ�bG�-��Z��s(�(4gO3 ��ũT#'���so��&���(m:m���F�h�!R�f�C�����6�f�E�yv qd�~x=�?�O�r�#���[�r �H�z^�Aޒ���Z�X�޷�?�%��g7���b۳Z!�:�������W��h�X���#]�Z��e��z�a�'��<���u_μ}�W2�g�~��`�ԮpqC��oN��e
a�{�f:��ͩT�=��+�i^+nD�ؕ�A̳��J>��c�r�yWe J÷Y�[�Q�<R�>=��ꏢ��}�qհ������*�B��G��m��R���e悜in)Q=c\���,�ig�&}ƀhx���]���~�����H��#��"#���[s���z��lD�k!�jS�Ȣ'�;oB����v������U��7(�0����sfշ�r�5�!�w/� +��qA�V�I�_F=K�+=CTF[Gh�E�W��L����<���&�s��=d�+#��4�#�f�yw��z:��t��XG�_7X�O��>���%�jJ}��5�'E��6Pᔰ�4U1,X�a0��F~���%
�g�$��	1S�a�����T�&G�U/�`rZ'��z����1�\���~�K?a�y�a��3�Di��?h*�z�U�&��h(Q ����*�1:�<		?_���p֏���%�����+߁n���Lk�E�P>s�Y�c��7A�<�2a�z���I�~'+��,÷y��ޅU�W�ä�T��g?݀�K |�=���$x��F��Y'����QV��xg�\�Ls�Zp��KV[�؉i+J��/f�l����{���}X�ݚ!���b�龎=�'�؉j1��Ւ��yEig��}��h�l@�fC��/�Z�]Ɠ ����E�T ���	`�d8.���Q'6�V��W,���͡@�/I����̀��pE5i����F��p�ŋHؒ$YS�8d�d�|Kx�w�+BO�Z�v�_�d^o�I�\O�����L�Z"{�S� 3��p�ɤ^w�L�۽�+�>�h>�^[3��~�d