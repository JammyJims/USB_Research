XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��OOm�q�5扒�J��X!�y�u��k>��|�����$*�P���$y�1�#����D�>��o�hF���X����c)�H��çθ�����o��rd�� ���؋O�׀�w���Z�?Y7n��0����Ɨr� �@��0-1�7
reG�#��~�s����`�`C��+7<��5Y�Z�DH�-�FF���W"�Y_���\�6	T��;,��,p���Ru��fm;V9����(��m�*O�Λ�xR�~��@.�(�yu�e�)TI^rC�d%4��$Q����)�Ì/�f���=��ipG62�\�fQX���4jn�{t��d�8x�2�\��>E
��lf�O��b���]>���]v^.1�.[��%�����Gѽ��PltZ�-R�sߠ������cԹ���9ٔ3`��%����y���| ��r���i���2ҩ��Hj{P@獽~4�m5�+!ɗ���ß��[�Ժu���b���xK��w&�R׭V0%%`��g���G�ڸ�a�e������8��rC�:1�q�z%�X�"�,°q�\z���������B'3;�6�O���BDPp<P�U��u��0����Zϣ�C߬��uɜ����K< ��*Ā!g_��"�ԙZ��gEi �*8�	)o/�~�d�.��Fg��8�����G����(1s��dF���~f����K�f	ɾ!����Э~��W�����D����¯+�?��T^���]mk-m��
g"XlxVHYEB    1cee     880T��䢆]U� a��fs؟m�;
�ZW��
�f-]�1�����=��J�
(w?ʸ g��=+))EY�9駀j(��������ʓ<'>'Cm�%ʊ�)���fisN�(�D>	ڟ�"gP{fq�k&�CO�¯���� �Q�dh+�\����l��:C=����(�Ul�M�=N�bg��j߰b��_�U�>���m=��b\}��gkVu�B'�8��B��KX��T��\�X0\4TZ���g��(�k��j#�`wW�?!2�8��8�t�&W��1u��j�mg:-j����
E�<N��/$ ���+� 
��3}� �e(�W;(�
�G��4�!��B.@_i�������]{�R���7kv��v��) ��UX#J��X�jڑ)��Y\�!T���
�cڶ�*Ô8|�7V�U�D����E'$"��m�g.b(#�Ĩ��6.S��8�����{2�{�n=.��KH8� k�y=����~�,�wʏ�D	TH�c�$���?_�����PJ�(�W�+��Y��1�UV�4�c��ю��O�2_i$#�I&�󄞔�-G|�m��tt5l��ޱX���}X��AKL6�
�i�n��AQ�FQ�����L;(��G>��֌u��p�<88L��?�!Ž�"#L_�D�w��W�ic���Bػ�@�]���.�M��Q�3Vs�\hQ]^�*G�ϙ�`YbyN��Uv�i~�)Է�خ?=��"�yY�?�e`��lt?A��k��J �|�+�W�*&�R{:C�mrԛ���'�:�u��+hs?`n2�v�J��c�>g2���G���MW������t����Z�R>I⏯tΣRM(#���k�0�ՠ�P�����O.{�k3aOȹ��q�Y�I(`�.�+|F�9�&����}��>Q�x���0懖�c9�
id��lA�-�SiP�FM���Ӧ@���;"��/P�|S`6�{c�5�!�4��]���Z���
Lp��2d����4��؆�ސ�!���qV-{�9�(��5D?%Fm_"���T�[�Q���"æʪb$E=DQK�iI8�j�{\eU��������d��3��}�5�/>�Cݽ.
yM�_�z�
UM�QU��/m�̤!�<o�@����W#�э��8n��y��@��t[��Ƌ4��'�t)���"�2�� 5X�od��˰��f&#>���Lh!������+���Ĕ@4v��n��aėӥ����:�~��\ e~}�aTq�6��:��b��O6���	k��?��(��y��xV��3*�7:��gfu*�EBas��Dv�$ %��f嵗��K���bkj|_|�G�_K��C�q��.�N�Xv�blH�٩�<���޹��H<[<i�:1_�Z��qOyJ!mK_�Z�ud%K�x��"B8q�/�%)R�C�8��+�/r���ֶf�gG��[F.��s������A�3�ͅq��������e���RdzO��Jmnx�S@����G�yi��� �v�s�#֎�����<W��n�52$7���W�v�< -X�/��mw{�`�Ypa%��;2T#e�9��Q9m]Wm�7��t��0��_��[�'\�]�rBUrj'�s��:�: �(�.^��ru��[�>)��=P�8=FF�lg$VN�[���G�j��?S]���<����^�Z�B����+<w;gXR��8,²[/%�(*pݝ#,�9i�5��ƨ�8���uN�yF�0;���܎�WR�M4�f#]����~yKX`"���=�Y����y��{�ǩ!�O/� ;�k��+ ������
� 0�VP��R�x���t�
s�8=�h؇İ�)���<�U�7BI�%�1�ѣ��L�zO��:)�?H*�/?��U�@]�|T��.�M���l���FMMw�����L�D��gکq�ܴ�ֵ%Sf��|�Qd����Ǒ��G	�H�N�y%�%nr$sT_���Ԓ�����ƐgҌ��_/h>6o#�����%\i##7��)X�DО�s6T�A�<9�Jh���E��H���$�x�^zԅ����ܥ�)am�왇�a�d$���,`a������T�I��K��|hw%��.,"$�6�{b��=�4�%H�'�J�����|+�F!:��%z