XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[�T(�\����C?�o���3x��}jE�'�<A)�(��	��O�;�����I����i���}�%��y���7 `=�|��L�]�r�{�*�qU�q��;\XF����%��B&X�&g8��.:�Ik����BZ��+QIyԾn���۾�v���v�e�$�ˮj���m�������5�^~��K���K��uJ�s�o�/�) �|�/.���,?n@��H�z\w��a�	���i���Eœ�)+!b�����$�r�v!/��I�jiN�/�C��~E�꺵��`��-���^�kL�Oo1�5�
�W���G�<c5#�����_7�~ fRⰫ\�e}a���ɿf��Uq*�x�F�a�9�OO����ٟ�Q�����D}��!X��o[����3q�zP��ud��~���DV�w��g����L8��x����c��[�~�cq�����k0��p;Qu��!�Όa~��>N�Ec+oX�8���*��%
����Ux�~((��!��7f8��\�?������6���d�������
U���K�j`�ׂ��@.<��4.��	fп��uVO*���޹~'#*����u@g���!5�R�Я[��"��He {R2��:�խ��OiK�DL�r2/9�<؉�I7e$t���)~+hWR��h)���X��/-�
��pY�Y��� q�M�8��Zk?)� �*F0��G�	U�kC��j��Hn���1��Yz��i;h����LXlxVHYEB    4c76    1340W܆�=}�Hi�X���ӟt��_vGH�K�g�7	�҅F�&�#~z��p}ڍUh!�{��lV�U�Iȏ�oE	j���t8�ي�+��q���?�����nR!cVG4/`e�޾ ��t�yr��q�9鄅���c����:�L��kC,UV.�F��p᝘���6���>�m�#�O4�����R��=�>�J/�`j���i!Zx]�2N�ȹW��,4]�;9�C��tǟ�q0��9�Ƞ��� }��ᴥE�
�[L<A,�[̯^��9��v��q^0g��'�G4�ɼD�����[��G�"�~����sJ�nn ��KmB�X-���|H���Ѭ��u��`�e��?2|Gw�:X������?+��I��y0T�9!����W��EmC�-�p|!u�-���,���C�0�|�Y�_Y�!�	/[�����_��a�F��wt�ί�w�%��R��!ZU�)O�iQ�n�%6{��M�ѿ��̦V���,4>��ᖴj�U|V��04����1y��A�K���EQ��2l��g�?r����t��Y��%�e�w��3X9ʮ�V��pb��K<�g�Y�LUR a�KӞ7��<la���$���T�+�.
��L��gM?�{_%�V}i��,6��}��T�v��!�ʈy{��>�
�ه�G��:�W�7����;r���HkR�h舰� -f~��H�l������TZ҆&þֲ����������r���gT�0;�}����4V�Hw�,������kI2����-][�#��k��f��iG38:�w�֧��%҆-����v�C1�1gt��Vf��`����q�������L���:{}�!ڪ�N(ٻ7	�@��VY�����)���C�/%�%�^	�Z+�$�l������2���?	I5��oVG�07����M("/�`�ɥ%�R��7�L��'�u	����|v�Oj�T��\� �|�,�����0�b�''jץ�l��g)��-�{lST��<��0������a����Ɠ�d��o޵��}��d��[�9~"-�bi���CZ�^[2���_�Xql]&���8+�I�(������N��	��G,�T[D�F95����k�Ī	A�iE�{Ȇ�v��F���T�"g�r=@E��䯸�t!_^M\	��TuOC$�����?�׼T<�i�'r5I���(<����<\���8б����ޢPv���L�F��JS�&m��
k���!�F�HKYޑ��!F��'ߵ|˺/!Z���b�j�"#�3O��|+��~��ƨ��Nq+��떸T�
+e�%<��~K�ye�1=/b� A�}�<��Ř�PWM��qO9�0�{n@M��m&��� Ģ�6} �6E�ZV����}�/n�N�i��f�����;�p��$�Kx"�n�AX��:|g�k�p2�r����fa��aFD!�#�|�����#��ŤH��$j����v��Jl����F'k����w�F`��i2����~aC�XcH��i�l	��i���cvFY�O9ˊwˡ����<r1�B���r��h6N(��Q�+q��W�i538f3�R�b'H/�O�?5A}�DP\�%xA�0��0�(��	`��3��Y2�,GTH�eRK�(!d�:��x<�iʄ�����74�����Z�a� ��{��#f�#�YE�ܳ㒕�h��3/���	%��D�6��\�(.Z��L�ϭ
�?��5
�!ښ��(���(������:`�9wZǜ�<���4�|uM��?���e�_�[�6��J��^����4���A[���cɫP�v.b�Jba�����?�a�Szi��5���Z@Xۢ�n�=ͪ]�`U>�Q��%9 �Bja��٧��v��EmC�M�r���H���|����ݥ�+0���
Y��/��&�f%�;����V��,�!4*������#�'v;k��v���S�Yn{�M�c���n{@�9̈Ͱ����B���z�>s�ٓ��w/�.�=��f]4�C'l9��"[����6jH���"mIp����焢[��[��Ӝ���nր>1�b�J�.���ݰ~���Z��E[�K��n�t]��֍-S6��٦L'�o�e���3�wou�x�a4Bj�P���	s���cJѥ��&�r�GL�)Y�p5�vӏ�!\+1i�w�ƫ5&��ԥvuUGq�iDq��*��XZY,�v�9�m#z71	�B-V	������z!}Ϲ�	=b^�耫�qC{�P+����<�~~��\$�PQ
�ģ� 3����~�Ɵ�g�5�\�%���[%V��$.���Z�I��'�{�B�����+�G3��#z��c��o%�P|�}r���:`8�u)ZW��-�Wܤ���^��JMB�
� Õb=bxr�Ү�?	�"{��}�JV��E�vdDj��Tr���l��n�a(=w�%-��!A8��ᤨ�HI|��p!$��)�cpx�Kˋ�Z�ʳ�#��X��m~)�r�WJa���9S�e�uɠ5MK�I3�*�����G~���(���A ���<Oa����7�!�7�6��ϙ����fKF�V�kx�;�S
���v�H̫�Ze IgY��C(�Km��e{�y�D�����ŵ��XE�ʸ�O��e�CqBɹ.�
��A���w���a�;�iA�nY7p�
J���E$��|E(�`c���1��@��#�v�xiDM7.�_b'4��$��Ɏ��J�Hf��K��e)�s���w1������'���x�>j�Wr HaQ=a±?�U�hl��=pM\���� }Rd��9�%lQk��^L�LV=e���^��ݻ0Vj9�[3�Y�u����2��S��r���3��Њ�Au���y�Y��, �������h~�%1ĳ�U���@Z�!��dx�������.<<��>�%�ޅh�G!KT՟E��gz�֐J3�#���"m�ͨ�	h�/�W�9v_#�l�6Qx��wqA�
_�iU�H��T�󫋈�̿"����S��HW�_�a���e�w<����Bs�w��`ԉ���h$���Q``��Ö����W5��*�CqW��zc.��
���x�k�C�<�s�!L:���f�\�喋Z"����\D�Vk����7���v�\b��z=�X;Tr��T ��Y�z3��o+I%�ָ���^d�����B<��"q�|�١~��	����i�%���s���:� ��̋K�m,�d�F��aj�gRkG�����6��4F6���i�糷�Cޗ�ƴ~}c�&CH/�u�W}��t6Z"j�Hr������N.���j��|eL��2��1�f����u_S��>PH���+a�]�c�/�B͂l�ތ?���_9yAa�<�S[�~�9G������
L:!yY��2�)� �� &���4P���%�3:8��F�����.P��]��A�Į������CxZR�Ia�0�U�o7�U�aq.ML+���� SqE��G+��RL�=��JTK~���>��%uϘ�g�f��L;e��B�߮��Eħ�`��������'����]՛5磦Gi����+}���m�L�S1i�y�4մ��!՟W���cjׯ�<�hW�����U����^�P��b�78�ŕ�EM�:�zXͼ�����[�M@«�5.���E1C*%��:���pahT�ؽR3�lC�gU7�������p��}�6<��1�Q;��?
0�W|ؿ�▧,��1}�{��Kx��������Ԇ��n(p��i���6=�0��VdMh<v<^�����=��Gxb���J�YDXTh�a�Q�28�PB����9�����V�#oӒ!�?�� iI�����P��'.Zޑ2����FY��Z�;����zn�`;s�X�J��j����i�u��U��"�� 'd9ژSl���*zqT��Vݮ�=�C�)a�F����3`��=-�<Y�+)ҽ�8�g�i�,�%�� ����p��!'�ߝiQ������/̹C�����Ґ�T���o�¥@�ȋ_��[��@����
Mn$�{x��#G�#:��4�qJ�Ϧ1f�I#�8�D�(��ܷ?dm��\ZTsHᘿq�K}�&r��ܪ�F�\��o1�f��:��WY��BgN�B�}��:U�;9�h>6AP=sP�K���緻���Nă�0�)��Z��zY�uiC}mc=���e�+��eS��
��E��>�AI�jM�C{��6�]�Tַ��<mA��6�{뛽���b���r'St���cL��}n�GVT�G���i�jX�VJ���q���y��4�10ʛJ�If��&���-�F��_\�;�3�Ư��X�ui�7�ry���ԙ�zM*Qg�F�$�j��5޷j���0z��u�>	���%�Acd�|@��M�A�}˿S��6p��t��${�v��pL+�m�sr9��Ke.kT%]`o��vK�p��c-�|�g��U���8�Ʃ����_����l]R����g��,څ�G6]�V����Y��vH����ٗHr��@6"��jS������S�t����#�rԄ��8?�Ğ z�h��.piDC}a0��O@�%!@�D�ڛ������Y��{��Q1��D	�6����o�/�� � nT����2�E�Я�)�G;f�a�*���'d(
�u.�N��u+�<�c}�E_�+>6g(Ĉ�u�v��W ��٤ �J�"�s⊂�-�������"�9Mu�I�=TV)߳ݫP���(���fc}.y2 ��S�pf~ʼ��XY�;N��`$��BR�+o~P�Gtފ���4�-