XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r?=�4����@��?[���0E	�.�"�Cf�Q��Ʃ�u|��`PV��#�-m���	Ǉ@N�W����Y�(Ă��<�h���O0�!�f_O�N��j�~3P��Ă������ �ҳ���D:;�joh��i��.����>��O/�]҈����}�e%�3y8���#L�1 ����%��cY�%�-�8��[�3�^/V<9X�d�8�*�҃�5Vp�v�Z���Q߉y����p��		c�Ž^�UN���wAg��q�� ��k�����ɚ�w�Ե�=vn�,��C0����T��V���2�M���<�'܀Rv廐��Ʉ�~<�u0+L3�^�O�L�t��qrT�fS�&�Di`ȑ�� ��Vt�������'�z~c �#��#9S+�wl�GQ������up�G�ޫ�n�M�`N����O�<���|5�A���I�MTn���['>3  [yJp�����|�v�=4j���T�tl> Q���\�j�(�Jz-�<�'7�G�O���|.�v�n���~���[�nV��K۹A�IM�J��W/�ݽ�]NT7����=m���xE��{�
�8�|�dN�S�*sN��s��d�*T����`���a��[r���̓`T�#h<J�t#�@wx�*=���D���F��H�v�������������`��7��L�"�Sr8�F�%��19���vK��H9{C�W�)f��������%�P���C|f@3��� Y?�/�]��Ӷ�XlxVHYEB    36c2     ec0'8�#�&$���K���/�I��deW��;�P!������+1W>��қ��,�4>��6�J]qDz�y\o��3|ׁk�ț�'D��[�ꠖz��JWb�����A��7�<�&��w���&b��B>	�W�@�L}��4�u+�I�f^4N��>\�A#�"}s����d���Njq`����>�YIT��$ψ�Z�I�ݠR���vެW���� �2y���
�kdrZ\:/�;]�x����7Ы��lrG�|،*�X/�|�8E�u*����o� =�?]�l�mXM�H��uij���ٓ�R��)�˻{�Cd4�a'����<h?�1)��((5	S4��#�n�שzĶ�)�|�sr�����N�)��%. ��*��5��)�n��K�Y��\5a��o���5��nH�p�i�ƾ/Qo0�G�����y�>�|xL���������m>�M$e������£Rb����Oo��9�"�YD�WF���N>3�(�����6�2�ћ�)ȵ��U4]7�Q��7��uS�7$���^+/-��&�q�/NdlV!�-"�0�U\���tA�d����D����� ["<k%�?A�V
�&s�5��J���S��MJh�wѿ��"�>�*�;�|ϫ�&��'U� ��;f,%���I�m̚.�4pP�N�W;�R�\{�]5��L�]����tSVaYfqX9��-Y��jN��ެ���E��z;?�Dc�z������&�+F䜇L���]�m�m"g�&���*v䷊���NP������R�$BS�1��Q����s}%�%��������wi>|�7���	�M��9�I���q2�k�n�p:����.��WO�l�a�=fP;��d|+���U��1���4
|=6�"��&QʾqU�{��a��T���$�3�a�k/)$Tr�e ���~�y�O�6Qd���QF��wy�,����ߡ��(}�N��c���E��քN������� �q�IQ�����p2~x̰�ܔ�����a�Ԃ�$�z���1@/_�(F�Ջ1��ѱ̄����#R]��5&�"M�uX�s�����tk,cC$`.�@]D�$��m͂�ϑJ[�dUb�����N���x^j�^��fhͱ�P��V�TsIpW��xs5&f굮&��
�:���-�v����u�ź[>o��
�p���� p�4�+KP��q�jn!�^7�N ��Ƃ���8�q\�+2et΀�������I@2����?軬o�R��>&�o�Y`l���Bn�5��L?@�%�D�Q_�ZrN�����[�;A�MVt��?q�DϨ�1ņZz�TPDF��/c�by�^�ɷ}�_�ȴĻ��DF/�Y�܊���s̸
�H~��yF��b�	�4���V:��:��m U'��R��y��y�KW�hؖ�����;	�$YH��J��R$��$�17��8�J�:�>�5f��CMӐ���F�5�{<�{m�x�`�z�q��.i�{�ϣ(�͌:�H�[�
��7��w��)�e�E�(��3�ڂǳ4�O�~X�E��w��s�W�\E�9䑨6(]�a��ͮ�P;<�q�|��0Hs�����|�-ŻR�%ɱR�����#":m�`T�̣�ЀP��(�Ҁ�p�p}���*��ޤ�@��_�*`�(�jEiw�0-��Q�ebR��ƙ�Xy|��hPYY"�`ɮu��{"��j ����VX��8M�*t�1�O�����4剖/+�`rg�؟s@]�~Rԕ���e4���ch��ḌE��T�Z�X$(|�胳���(�ӕ�������O��He:�����P�5�/C��Ẍ;��9��*>Dk
/�,��(��0M��^2�t��q�洃皎�\kc�|Ń�怴�l�@��i砆V���G�L{0��&"��B�r�*ͩ���.�����i��L�ix�}�,�E,5-%�B�X+��'�آ:���$�<���s08QB�gm��*m��e�.$-}ЀjX4��0��9�^:z�ˆh��/BH�%�}P7L�q 9�����o�u�	��I4qG��g��!�:��@N�b��Ð<���?ղ������IKYỹ��T-8��F��!Z��=�S���V�ͧ�c�*�Tғ>΃����8��*� <GY�hA@�.�`E?�?FX��&$�X�!�q�#,u*l>�J8�4V�?	���(Y5��J2�u���UG��͓�>���l���>�ku^y�.E�$iՔ��Ɖ�â�V�%�xi
�H�X���m�~+"�4Α+�H��Ibc6a�!j�=V�����
#G�;�HA������G2� ��_l�
�?�)>K�Y2w��%�E !�O7a���P�(n�)�ƌ帠��8�G&��b>��Y��%��]XL-gyh����Zw��0_����H���b(�W���K6���W�`�L��i@��q�`�����?H�E��af:��H�~�{�B*e� �FM2�����S��a�������źѤ6���Ύ��$0!a���P���Q��ksIA�xn�͝�t:�k�Y>S>ေ�G�h��?	'�'c� 5)-M�H.\����I����c3ct�w-�qТ��7d�SV�:�lڻ���ͿPdU� �;_;��p�S��0�y#�b��[VЬ���'�^t){f�F��W�=���qdb��� ��ʨz�Pp��8������-E.�y�b��2�������u�
Ϣ��d�i剮��}H��f��,0Tp�Au�0�u�O4�S���F�a�����=٢�\k�ځ��t��_@v
��oV��N;4.���Ip�k1�k�OX��
��P�R�{��%jm�"�U(�I:.���*x�3�}NR�&���ٟ2ܚG��:d�ܴ��9��D������5fֈ���S36��P���/�/��0cF�:@�%����N��a��m(C��k=wM)�+ÞlhPM U�US�
�VA��?��!~
�\�&F*�OV���"C��� �����O�ױtienOj0d� ׁo�"܁�Ư]���s�:Hyn��2��6|�t��Of�]͖"[�C�_G����tC�����̜���x�m ԉ|�{��iJ�yio�nae#�r�v������с�\�@�sU��xci����l@�����(�զ�9���i�����������%?E#[�y��v*}]N��� ���;	�@���Jvrn�+˓̜�ps��[@b�w�=���Na / �z�gpa
��1���]�uf��¯���Y�=�g��ý�������1��Ґ\a��U/�J�;�|��ř��\` ��F�d���$��fn	͉@j5ImQ�u����/~��G�6�t�"��X��A(P�����4<���B��`��BPS:���'ſ
�ZȀ��b	��$z7��	�GI�K�"�q�j'�G}�Mȃ=������䰼��UL�C�E�O�+Ik���W�!�`�,��j��.L�)�D�%uj˺��ʳ����9�8+���z7v��Km�)������Y�f��J���A4� �.���+V��i�eX7#��3Ìu^�<��v���Q)$��5��d�ht��E��&�_U�(�$X��'�ё+6�ѳ������A����пT���م��0��dlA�q)F.����q��G���@��#�.�X>