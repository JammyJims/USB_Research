XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y���x3��E�_k,�y��A�(��6��������x�j�М~��t�=�R�@N��l/�&�f�����L�W�s7��çG�D����bIzw�$�6�)��,�%�F���e�o��=������C�RA ���� �jDI�6��(���2���ǩ�9q����n�jX8#�Ɣ#�a��	��V��R�����'ӽ@S#{�����;' �N"�gP�"b(/@S��d�j�g�{nI�Ly���i�`.��0�;m��o���A�QD"VРR��GZ���P���Kg���rq���������"�F��A��'PY��j~w4��lik��F�^^�y����g�� PUS���Cm'�N��Am����������F�׀����ޥ�g��oc��%���(��B�a��ę����r��1ck�*�
TO��/����l�+��FS�;2��0�Ĝ9�t��&n��`�{����aL���v��{��$�e��b�v;����� ����#u��$�Nw�U|���NZ���M��^tfT���cs^��f�aE��{Y�E����Ò�������Ƨ(���ӋUMN���iJJ5O9Q����+�V��"2n�LIy�ro,��p�Y�����*l��ʃD�n}��>{%t0�stW�:"�[�9�����̓h����K�!96>���2��O���g��r�(�F��SaP����-J!d��/R__�����+f{7��Fl�;´w���g%�e��{�]C�3l�zXlxVHYEB    2b5f     c50��@)�Q
v4���n�j1ȼd���^��4/�Ԏ��0���4�P_! t8�KZ~�ٴ�P=��ֲj
M��ɝ�4uJN�G��t!*�PB��[��q�s�ڽP���;k��O*Xp����W=���C/v�+T�����g��J2�^�p!?�����+��W��M},�_PjP�*�|�&r7�T6����팛��AK/�O����� l��ȸM���J�Q:ɔ���$����
��'ˤ6� c�x��|����!J�h������~�$�6K��m�����~6�~��7���*����u��C+���v����z���z�*(��èw����R��(_��QpT����t�{�X-+�j���~��w�LX-�6ytq�JFF��vz��7ّY��`�����Ab��	���ed6�1"�rH*��*3�Z�, e��h*��I䎲/^��Ҭ�(�v�3a,�5ĥo��!�g�G)|�Ӂ+SOr���Lv	
5E�,I�Zf��8]�{ᗕ� ��ec��ҥ�y�[�+�T��� G�|����B|����T�~x��������4ە����$���qAR�W��fK��O�õCF��E�� �3���%��
|���Д6nx?+��*��@h��ݧ"eQ�#�d!cb�Q���2�:{9���w����W�J�"�ץj�7�;5tj`y�>F��iE������HeF��6ڛn�w˝{L�oo�r�3� ���knЭ̓�cxAE�x�5��+6j4�oxp��5�n~�̉ϊ�$�%72q�ӹ�^P�j�;XR)����X�J��s�ӆO�ּ(�7��|D�22�n*��f����~{__�/q��^x�1U���9L����1�T�i&�'ιə�������Ѕ1%�!;OJ��֞��?h�,Ǐ��0)�����эE�4�I�����I�!\�=�l��g�O�H��Sw~���Q��ޖ6j!D�cB�ڂ�pZ8'N���_Kf��� hA��H'����y�$���M�|�I��ł�x~�����}s�}���b��Cߤ��wִ�}�u��.I��ē�V�vo�2N��D��q}����I�E�71��	L����=fh�5��F�ɤ�W���NC�K���;8BJiV��c���������oO�%ըv�pa3 �͓o��(аj��}�*Mf�Əxβ%�T�l]����hx.�W��}��?�Z�,)�CjI�� #�`\��&���7�'-fR�����Y ָ4=�,o���4�Gw������ׄ���+oe;1�~�����N���_��PI\����!���C_�"�g�P���U�5@8һQY�`o��ԝNg�(�h�[QA5�+h4�m����߉x�)i�;���M�/��o�=��l�_�<���<�,xGzGW���a�z��f��=k�V��W�@���|�zm��?�9bc�	=93M��D#q��ȦS�ؓ�s����P��s�ϡ� `��F��eԵ��ٚs���ݶ&6�?q�.0\8Rr��~�}����#��O֢�.��|~ψ����:L7�F&��f�G��e�Q��f7�U:�VS��a���f0��r�%�"��:a{a�4m/�<x�4��G�\K��E�8��S���,�̚Z����]�4�ݼ�v�c&D8^�Бt�O��T�����e~�+�޼��v��-\�܅U�f�訷釰ht�+��u��l�����@���u���se:���g��q4�H=�ioqՁ��Yq�[$h���Z nL�K�Jl.��3�o��(�Ng2�y,��{v����U�~�#��4���ҝj�0r�����ц�$%nMw{ȋ����8-��z����Bt�@��g�����o��x`��Be̽��K�����Т�{���D�7[�3N�HK�����|�Q"{����b�(V)p����{21�fMu�Ө0�����q�7S��tX���Ч��0!E"�u�Z��Z��q�${s�VoL6ѥ�����x�҉\$x��=�9)c0z,��ղ9�e��H�B�ue_·��I��;��o�m�Z�A(���-�9OA�(=��a9��vk!�l2u<j��D��m
���dZN�m���Qe����2��C���.��K&��Ɨ�JQ|�IU��0��"� �`�G�����n+�O�He���UA]�"�UO6��`Yr@T����!��A��<_�Ϥ��HnAH���*���x� �KyBCs�l��Pc������e��5A� >cB�sy]�,嚷�_���EV�O�``�<�T�cw���ϒ/�����V_`U�����⿃nz`x2���[�s��!��0��~}ӎ2N��z�>��p��r����:����~$|�q��R��p�zw�B�9,����û��W����2�nk���h�EP<�Ut��X�_�K�"�u �BB��G�U��b�k�)�mECE�˾zPV��ޝ����&��8�q��
�u�0�~��1ɰjZ(��hd��~������Y��:�O��zA����D�H������Y�����8�y�����W�?�>��R ��^u��͛F��ʛ兟<%G�����t���2P.����"O��cK���Rj��&>ۆ��JD�!��K��ڞ���ak(���[����X��nɃ����Ж���?�h*�=՚�G7��JX�
���T\�^�/�-dm��`ת�Zz�������C�{c4��,��H���j�O�Sm1�_�A�'�
�O���F�`R�0��ܓ����N���t)Ą��t�����TLk�y�K`SN�bq����ex7��s�'�Cw�L��?4u��.��x��L��E,�ʧ�#�k_���yu��7�R�lib�W��0U�K|>C=e�iK��^oX�xU^�Ҁl`��:��� �<���Vs�5^:%H��{�&R o�q�*wb�;"i�7H���6��d��b?d �`7 �s3@5�2;��vfɚ%���ܹ�]��v<�}�%hv�IZq�_/e+�$|����jⷴ����q�aA��K����