XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������l|�����5a��l�gM_����$-��Z<q�.:l�,���(-�:�3�i\��1P�pG�MiD�FN��P�eC$9Ԕy���c�w��������30������-%�2]s����Nz8T>U$S��7v{x
7I��4V�$J���]6���d�Bq�gR��Y��
3��Nm[T�vF��)~��P �2 f�2{���B�0����؍� �*v��� ����zú�Yz�":���o�ۛ�woF�D��T��*�Ik��'�%%�`S�{�ε_��Lb-�����+�x�KQ��j�F@��̄R7��'XZ��\ʩ���w$�䍮;��L�f3��
�(':I\\�0�J�J�m����j����g+���U���ڌ�{�����!m�6�m_~��3�˛"���FY�1,�"?�P�ڒ5I ��X�땠�&c���31�a1]��Kq�#���]ڠ!�j�i��h��B�0������,�5�����ǧ�BI5g�E]9	Q�rl� �X�*���q%�g(�F���S��ԅ(SAv��a�_��8��+�[���	����Jsnf�Ӏk���s�e�r���p�:���T2�s�V�_�W�t-%�%~J�ǌe9��dȜXمm�t0��bK۾\0!���ĺ�z?�.���H�-.�Te�Z�B+�?�6D�-�qmQmN���7L[?�7[�����WX�Z]��sί%=�ᓬ_��o9�1A̬n$�XlxVHYEB     d62     660�F.B��h�r-��̎�|3�V9�;��,���\mǨ��.1�'/H�F�@?/��᝕�D_�3�+'p�χ	��{y[�"D��M�Q�˒�oؕ�N�
g~v��5A��	"�'�w�S��;.��RP��P���<�MVk�h3C��.Y��lܖ�N��K3�N/&\�ȫ�C��)P������:!����c:�7��(p�l�Xľj��0U��6ψ�����s�%f�b�K�*��ks�M~к�D�"nО���\��Hp ��A��O͸���ߞr;�Z�"?�l n'��8�crǗG���1���VMbh���!b��?q��* �p����u�@���۫�!�C�UV3uI��鶠�,FS�g����T�n]��jXO�+����Ma/��Q�uT4)� �o�zhw{8�p�*�ܻ�`T[���l�%BXK�m��* ���VM�C򺔏T!1�{��k_.�h�k�[���t���?�:�19fRFoz7��%��N:T��Z��}���� �m�KAYʐ<�(�k�џ(M#�H
�n,�Hi��'�)(t��Uui�a����V�7܁ɁKS�G��#O`�m����~,دBw�7H�G1�o�X�|'	��|���~�<�����=�"0ya�5��E���]��L�Ȳ�W$�)�&e��ve*���'�� 
cL��B�z��e
���ۙ�?�21PV��P7���
�� �y-x!��٪�L�q��eYp�����GqtB�i2kGGu2�`^
�E����RY��,�K���NQq�,zL��Pt:θ&��#���j���fj=�!oF�����������r�Cp�)�E�Ou�i�Mq��@ ����+x��8�~��:v�Υm毒�"��"�4�t�}�v��,��d�<�~q�S9��j3�QY/	��.����lI}�
Ħ>a�ؤ���]J-	��$���]����$��m�U`��p��x�x��xO��>�����/?� ����qf���<�;����,N7�S���O�ʻO P�-�@�m�U.0�Ƈ	�I��as��M�j��
����z_�Xs�(�y{~���U�7�X1�w=N�4a�a��T��{�.2�}�~!7s'�h _��j@"ׂ�z�p�ُ�o������]��������!A����4Ou>�뒯��}:�K�T����x��3i��P�Q����@�{ [�x%�D��������΅��to��ޝ��Ey:Kh��rS+r�4-�� '#BPT��?��=���	4���`��e��ݫ�M��T�!��R�yQD���l��@f�^Z'|r&Ø��U��J)��П:S��sk��I[Wv�2u���A�ao��d����>��(��o��2��|�{��������;& �(��}i������uL&f�n�8��N�30�$����Xփ�p�@����i@sb��7y���p��A��ҿ[�6�L������0rg�h̍s*U6���7���Po�P��g_."��t��F�U�(�1*���!�j��R�����U�dk��0�^جo`�C����+
��W�QM2�}E���D�^)�
eEMY�=g�]�Tu��s��4*�