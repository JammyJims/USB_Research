XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����P��N=���ۖh*ĴxRe�c�!��r�c|��|R���k��s&ԦA��z1�-��
I�Lh��h/5+5�V%~�VV&�	�[�}٠�s[�Q���t��G�Y�,�Qű�C�:[�����2�i�F���$���E|?��f۩1�l뭎N�C�:��31B��A�5֐GpGꆚߺհ7Mg����a	i�x�W�'�q�w�?�1���w�4�Sݷ?@E���5ض�]�3��R8ǀ�W�A��a�S�8��'�َ�)�6%�R`�h(z �$��7�zs��=8O�,��Es@}�<�X]�7��-b:��ۥ ~L�2��9s��\�en߼�����3�\6�of��j��~�����1�1Zŧ��h��F��^e��hl���S�ߞH��O�`
���[2�[oNx+��꦳�ߴ\����l5��Z�A�$ֹbq⫖`��S��q��4����(�a*Z��)����'UC$s�÷�,E��]�o�� 0� �I����%3wԼ��;d������m]ڮ:�R~~�yq�@�h�G��'������}�y�vz��<>_���y��M"��&[]�_
��|"�̈́�(���T1љ)ZxM�n�����L�bi��|��C�\�}R�vv5��l�:hN
e� �憐�`�8���֦��X~�΅}�-�NۀRIX��j��`\��A��v�O��~@���j���U=*w��[e�����q����d�n�ܓc����W�q�	������uXlxVHYEB    42d6    13d0Reھ�������<ރ�Ve�J���*C�3cQ��m��#a�ﱉl�,s�ީ�ቓ*M�- L��Q�~�`k�d��[��eZV��Dl��ۺ3S�3�j���K9����_�����!�D���?~��C3�W����G�zH^�gt�%��*��.���^M<zB���~����;i����Ф_�i$+1�vWQ�;�a����0U���Y驦����&��7mkW5.�m�v���^���¾�7�P�g��.G��
&;��?<g�\��)�fHB���$�w�&�¬n�� k��aY� �i�f�����s���/�D9�͸�TN�TV�ǥ2 F���B���w���ALV=�Wg+�Z�ǀ�G�朗lx��W|�U���I��d*u ��ACN�X-8��ig�Ŷ�\ɂE�����OR��$ p�֟���
������5]�U�Vl(i���8?���zK��q�^C��kS���o� %2S��Q�Zr���&p%��I���*#�L�	��P*�5�ld��}�G�������"���s��\��'{�$���UGvs�uWO�QJk���� 	�Ҵ��veE!Í�U�@`\>KJJ�m�ݵ��(=�Gj�nU2�gK}G�6S��9�@�X<�0�Q�}��+�h"�.&dY�M_�Ճd��c,��L�ת,�q�4d����(�U~�)��N�N-Dl��ll0`��!w�RlGbT��=G��<2j����fpW3wڹ0�:�1̾,���m�Q(x4�vB��Ͻ�I�[q�����H*���kt!��$t��i		G���o�s�ʂ%O��V�{i�d��>�ܪ(M��X���M��
=��\Oމv���_$�;�ЖZI�U'[�ok)<�܌����9����U�P�� 	E���k*����O��@yx�R��sZ���-�[�k��te�야�ٟe�!Dq�-� ���k�m�72�!R$
��RzQɡ��j�6j�||S�QP���
�6N4ƞ�'��gl���0�hҷe�%C��J�$n��]S)l���T|��)�'"yMv�(ô���MMy��kb�a}F�.+ڌ9 �d��Â��1��CZ�7.ʆ!���8�^@�	�0QS̖b���E�'��*dTJێ�RM�hJ�{ˮ���w�b�-}���_�c����-
`ʽ��0�3���J�r~����~���u���0�f�EE�ރ��Ǧ�%�S�WDag���;�Rρ�-̜*z6�ؠO��
O�Y!�i�� %���� �e�= _�x�1���]�o@S�޴<ө�'��XD���;Di���N|�r����������>EK�]�`�R\ҽݨ ������Tc'�+�'3��H��7XkdzjyȐ��j;o��8��3��6c�����4��� =�����%&_I8!�1K�a������y;���F��46f�C*~��*v�+���S��2��_��G)3B�M�)�;/���˸B�GhP�]��#��Ŀ���9inC��˱�5�&�/�Z�g���j��%z�,���}HR���� � %@�#��#�ٯ���Ĕ�rj孂S����4P����TY�uj�pBb/��z���h8�����I�=���ԅv��>bj�A4���,H$���;�f��S��كlQ���	L�f�&���� eQ�
��6��2w�fMK��?��^aکW��:V��ȭ��Y��[�=��{fM���������&�~Ua�9����r����=H$�'�tw\��kv�c˘����-�l�Q�)����Ӵ1���D{��jRt�$��kq����"��ш���&<�RX�E��ElCKa� �j�q�iw��d\&#���H��m�K�g�Q3�d*���ۇ��D&�Y�X&�7K=tD�?��x�ℰ�nȄ���`�7�N/U�^��<]&/��1�q|�/j}Q���#�6����%L�`��uqm��\��ѱ`��Gqy���x����R�,
9@i:�V&��{�#�uT���������P�&E�3?[��n�d��}��z��5�ͥ���w��d.Q�$T��1��tI�I�9.��0�0p3�63����k�Fj��o��0b�$�^ �sX��%��Xڮ'�MB����Fp-_��򲶍(rn��3�/߆��v/�T|.P�UVU��_n��X�L��	-tB��{����kLeOFC3�l��vӖ~�F��~�9�@gn�KI.���쑌��L1�ʙ�菗�lv�2�a��fUY�*;��@bC��Y=�>p��b#��g������}ϼӮ�eDq�*�ߝ+���)����M�I"C��Vؗ@�z��~x8�&06�r�n>�Ѥ<Ea�̠��T�Gڄ�d��t�OQۨdHo�}oͯ�*� ug�̦�
��S�g������L_$�1-�S>�IH�� ��0�@ia���Y#�hu�����V�JMe���{9m]A�^?�H������p{ys�k��3�'j����R�?��Ꝕ;��;�1�Ńʳ)���d_������'�у!���F)rvq�6���t5�Px����-	1B*�0׈�~��#`N��?�=��ص��%R(t9K��U��w�<�U�T+��@5��iSuFf��h�.�Q��KP�n��] ��$MIp��Àţ�!�pE��b�;`v���yU�P�MfM>}���gK���Ds�h���t�C��u�@" ;��<��i�P�$�Q�eݢ�w,�"�$W���Y	��zғ@K�կ�!��4�,??�%�lr��'���!�]�y���?s�l.;�vw�����Sj���{���0��&fԋ�@�*b�$so�`Z&D6YbףsvJ�J�n�p�z���0#�l�(�X�6Ml@iC�fU0��DڎuHl�[=8|$�*�$�_ɠ��^��]G��)@&cN<��e��)v����:u�8O��A�x\G�<8�9�i�����u�F��]bB�9Z0�	��(�rgV�$�'u���-�]�*�]�EB���0@�l��T�e ��\��&��"2� O�/���<g�[%���붠 Q	���]��߱���F4�����I�'tb�1J��:b�Bj\��'}�D�I���^��
��_���',����	�+d;�z>0�B�w#U���g�B�!HB��o�@#W!7�t�S�4y� �X�^�Ou�A3�z��G��y��ֿYh�"��Q�}�s[�\�9
=������n�`4�Z�B���@bD4���������%n�/>88�3i�9-`]���<ze�W$压JCX14��GM���QϬ�_����~�1��aJ|u��8����l��W���1t�|F��ߒ*G�z�E�G�"��u���f.,d@��Z)yTNX�����/F@�������Θ�Dy4`ϼU|3t6��j֮-q�T����&B�9.��ܱKFpeӇ9΀c�t���H�T}Fǔ~ǵ��O���K'����HAѶ�Ɂ�KL����ƨ���lY�3Ir>y2^�q�"��� �p�m�?!������6:�'0Kŵo2P8�.�%��y�R���3퐫%�ox��^�+Mq��_��m�[Zz1�u��t4:2����{:�F�W�j3��r�]
���x���"��$\�W���V��w	���b��l#��V�-��:�i���2+�\<G�	���T�6�rQ��o
�@�zN�9FN#Բf>__�/6�U�V�S �3��ߕh��67��4�N�� 7׆�izE���`w}R/G�I�&'jo���e.Q���3���_f��{�#�/rQ
`�G��,>7\�q�ivg�Z��)L�'*`�s��4�O�֕��H*�m���7A5�W��ĻÛ���ARѨx����E�@��FѼ����D�n���Q��q]
�g8�Cd�S��HxC�Gb���T�A�۳��)��?�8�0��T\7?�2�������u����B%A�G�Gɉ[�k�k��f�n�����P��e`o��5H�Q�I]�k�g�n��%��#I��"O�M�.����)S\���������#ZR��91���^��cGA �A� <q3�OꬨF�[W�jX�:r�ϥ]�I��%��P7%A�N���N� 4�����:J�@��U,�a�R��ߝX�n�l�~I��՚�<%��N��<�6�-l��Re��|-�$��5����]��/���s#]��Ml��M�3s���q%�6��U��y�+;�~���A!w�����R۝�包����U=W��t�e��)�}��.Zw�J��J�����[�7����n�:R�U�`�( ��$F�bCSs��(�'5�0�������2��c+";ɛl�i�4���	��"^03z�ʶ'e� �C�~�������� ��p%�QL���	� ���H����WO�	�R��o����Bhɟ*�N��)�� �* "I����Sa���tpvtΡ��������G�$�<#yGl	;�a[�N���aH���v�M6�O�B9�8'{/�XD�?ouJNS�3}\����s]ݧ�/0�Yp�!�g,�T���|B�.��.B�i�l�TG:BR���z�s_�mV�V��c�Ǫ�P�/B~�g�dZ�z�/#��*�l��j�<��lG7��i9�:��6�Y�"���RU���1��EO+�z�,���p�+Zp��s�©]d���N�6׌De%Z�֨�Kh)(ue�X��!����P��Z���g�fӄѧ8X�Z	�G�D-�]�Ά�/ۓ�����㤄s�6��B<��yp� ��p}��)��~�mTӑ�6=9�p������d�^Ǥ�$�p��R����Љ�^��`����Yy��� 2�߼!uNIN����u��ơ�'uP��?�(�b�)����?m����������[S����ɩ��5n�%Zzh0=T�{�i����!����UC�п%�?O�H��aw��C��� ���+2����X��F&�1������