XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ȼ{5��/��*�R!�B(<���6����Τ����:�V~�\2D"��?�w�����j�=E�S+5騥����u�_�J���S���a��O8y�R8R�tà�^>�&���Ϩ'�8�+��Ϟ�R�sK�XsZc�C�\Z/'�]@��7�Ir�}Jnݼkn�n��h�!N2Oĵ&@���v��!�ܼV���t�(�eY�|gV>�x%f�	+��QiFA���p>����y|1	;4m��N�}C?�
>|�[Ǳ."	)F� ��,��D�"��gK�L���UN�y��2*��x�EM������������������[c=�� ��ڈ�|�6��*���)��Rc���#n�he=Z�"��IV]�=3e�&�̌���Q�}�(+qK�$?L	EY�цn;f5�f��<y� Y.�>t��s8����Ar���X��?H�㡞�|$tmj�ɅBg����Ɣ���^���/zYf��vY Q�0X7��u�����7��:ȁ����}���G#9T��}w<K�U��$��XW�Jj����|)����f�m�(B$����bX���}�_��c'�
.Qy²<���m |7`5Y����47����i?id@dCPHNS��gST�.c�t߰�T����d}"w~�@ҫ���]B.��lbƒ�����b�̀����'3֗�����KzvwuH�!>i0}��$i���4	���3�$�ך�R�6Z֯=x.F���r��;3���u��VG��Ĺ�t��XlxVHYEB    30c2     e30`O�z3�۠�I�����^��9�����y��E�^�)4m���U��K�u���w��	X�0�\��RMR؎��*�ۈ��A,�$851����ús�M���HnK*�|ktE��>�i��ސ��8�
8빟�����O��EZ�t�k��˸��(�3�R��'t,#>!>3�C��D�7Ы�S�7�	G(Wٞj��B>~S�����hu�����`�Љ�����vL#������/� ��
2H(�:��������賧
�  d��+�m!A�|�ּ%�(��*��[0װliwKR�C��>=��7X>Hz��4�lhU���*)��ۻ?��P���I��#"@q?��ͷL���H���ᐔ�HTz�b�}0�d�_h��R&�����ӌ�i����21sz�����r%5�v|5�*�ŕ�f8�i�.H��s�ŜƳ�QnȘy�_#2�"`���+�Pe���(p���3�֨ۮ�e&F�A�1%%�8*x[A_�t�e��/t�"�'��d�2��Y�Q��]@d ~>�`�����wK_
�Io���<������F!�)�K�X����u�k�8�+.*����Q����v+r��顜���"o�z6�j+g�O���Ǯ��)���6 �nY�s�����"Y"��al� �ZA�h�X.z� �i::�΀!W|2������s�sb�gy+gT-�k�PV�|^��a��M�鑆"}/0�Ww�Rq��� ��h�'�>ô�Є]DN��
���s��ԙ��y2��o��px��6�� ce�q.Xd��.���	��nq��Y�Y�:6%� �<k$f�N����nɑs���� I�G����Nu��*jN3\7���U��kO�==������g�*�}�!�=�h�D�%���D9%�7/�Ś��L�w2a��zʁ�Y�sVBsT5ϩaT>�B��l#vI�-3���V�)��U;W�͹���VEյaƜxO��mǇ�7���C����<�MSrTo��h�rqRZ֙"G�5�\���3a��i��h(j/�O�rB7�p���,���v��;9HSG�?������r���γ|�K��h�[���	�����#󉉌�G�l�MrMrڅ���0?D�PAFW}��¢��7:`C����)̍]�Z���kkLM._�m�� ҲU#�>� �_��CH�]�<�!��:���W�p'�%��	��PZ�K;p!����/uE��9�b�}��&'�V,R�j������]�����Ք��L���0�T\E6��H	M2y,�~�
	 _��o���f`Ks�ғD�+tyq�,Ċ�?R���P��iA.`�(��kY����G#-�1�	�4�T��w���n85��!�r'�bٯ5g�Y��Ƕ㻎n�K�q�
r�J�z�
qecG�l�_�������V��<Q g43�<� �-���H�d�g��6�)��?1�#�����݋�&)�tHD�

C���d��ZY����{-HVE��`e�6dS����2�&\ jD�PU5K	���c�^fn��q�TD���W�=����>]q��3Sc�0��S�w�f\ ����8\g�@��^�~�Ƈ���8O�l{�-"d��U��s/�ߍߩ�^��TQ��L906˫]c��)mL�NQJ�j!�I��z��o�Qh���cKX����3Y
S�a�	�O��3G�c������d�sw�"�CV�("	Ӭb�R��zب�Z�����������}���j�� ��{N���J�Xݽ�f����w�
{_�Ǟ߫��,|?�6�@n� ����[�"ڿ�
����֭��KUe�Ҋ�1s47i�<�j{�A�!m�,|%d[�����v1q�����w��5$�I)��:����<��#����� 6�&�9<�(ܛ?a�]�:��S�Vֆd�$����u��|b��@��8Z@j�f��6H_�����F��_"q�,� ����~/�tJG�k؍�d0�<&�4g3X���ŉ�����0/���m2R�9y\x��N&j5@y@(�jfEP�!u��_;��� �}�^�ZR84�H���U2�&h��������m�WmPd�;?u�����,OOP���+J/����-�Y��ﳜ&��i��|�ix�N�g)�fR7��02���F�!&�"i|��a�m��V����`����N�<ם�\v����j�A�+ZH�����X.#�z4^�cR^a���B�l��"�	��I����6�ʹ){n�]'��,� fY�Mu�V��C���r����.i�#�-� q5�[3�����S�pp��}��ҩ�����ZFUE��':���.���uǒ��b��z�!芕2����O��܂`�%YvӍu����u�l��E���z��t�&ѥ��鴀�f3���Q��$���G��)yllL[��st��%&�|�2�Yzk⑙�b��vM����ՙA_�\H��	�R1���X�[וU�׏̧�~����������xf�(���s�%H�WA%̧�]_���k��?9lg-q�F�UA���B	�|Fp��IA%��`R�����KB):ؤ��c�#0G��U��ߝ�@����ƈ32�����vگ��#�Z�m�yp�=�'�Py|�5v�H�yuD\�b��h�D7�Yb�T�k��.�
N'��|����ʑ�����s�s���� ��x]�8���q'�1�N���l�]���6�8��Je������'�G����H��E�l��q\�26�QT:ze8KZ�q.�P���HVIP 6�u����_�7K�ؠ�S��mOȍ�g�Q3�^��|^G9A��X˥�q@u������2X��~�]�r:E=9^Ŀ��=��)�J�~�V>��MН��Rgm���������P:
�Ha���'b�R�լ�B^����`i��,:�%���x��r��y>��QP�D	B&�/�v* �rea=$��K����=H��*�Z��C4�ʛ�����VI�'�t(����/9�je`��	`���5�/��rrϼy�:t��.�E��a!�7�j�t*���꒗�7ud�m�*��5���I��/��[%V���(�ݨz���4R��NbxbU���b̐ごRS���~��n�V���RR.;F�x}�!����c� ��P�z6�ij�a'���g55-�VqS��n�!���X�VDG��E�(�Xjcq�=����b��~��2�D�K�;��AsiZsߍ�aj��wT���OH�`�����:*�֪�/n�@}(W���!�A�Ɵ�{23oqc:�K?�I7����7�X�O��H�j4�6�&YE)�_�\�f�{�Kk�*�Є�SO��`=͗O������fN��ԟuOAB���4)�R �<9���oV�/����)�\O-��HR�j U8���Wnu��d�g$�B�,�Xr�[f0�iG�,�\���}��0�]��jΆ�9`BUh�V�;��S�����I?8� ���b'A"�c�1�?��r�2_�+��3�V�;,K��S�y�Vϣe�z(