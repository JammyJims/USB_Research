XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\����!$k��rP�#6�+�Lѽ���|�8� ^6� p�#�M�L#\H�ߍ�LQ���S1�7Y8�}4?c!g$�X5� �
����HgY)eAѴ��������aGGR�sg1�I�>�Ʃ Σ.��oV܁L�Ǒ �nMF�gj���R5��`X"%^ �{b6(��e]p����}��/
N��Ӧ��/�$0��Yf�bEu�R�m��8�0&�-�3��"�[Ko7���=~rlY����D�=�����}�U�l��5���i�La���n�`+�'\�y�����:9{��z�q�p�g��+���!�����Pt���p���/wq�[�J%�e-�y{���>5���s+���'�&|4�tz�$�|h��ʟ���u8��^q�ñE�
>u8l� �0�1l�\�j� S��C�	5kh5m�ٿї�"i����rz��v�be��f�k�h���*�x}�Ԍ��%�8(�{�d��k��.gJi�Yg��>��	�@N&�����ѷ�=��g*�B���� �c��J	�9���D�g�صa~H(��Ֆ\uг�,��
� a�di�د�n���F8���ˌ���������&�u�``���.j��݂J����� TMoN�0ڝ�x�t�
곸���_�xm�bЌśj��^��I���$��R*�3�2�i�`]�uo��t�-��vxNĖJD��8�7N��z�7��È�<"��b�o��FL+8�����໣��XlxVHYEB    fa00    2ff0���Ўπ�B������b�6�}%��L�����$q*��L�Oڸ���Q0�s�?����G��&w�}�v�!@3�zdl}�q�����9�a�$��d]
����.��*-��Q^�p�����8N�8��h��>t3,�ϴ�`���:©����0��z�ش?�ಗNꈜ���Ƅ��վ7'�Kmd~c��?��I=)�yxٜ0N�v5��R��m~�r�V�
P..[L�SA�\0��ù3E��
@k���52yvW'�V���$��t���Rw�`�x;7�pYֳ�����U1�A�w3^��e�o����?�Y�58���%9�eڭ*k-Y���߭E���T�Lm��I��������8R
�j
K��dE/_.QV��h�����F��`A=��-���O�+a��S2WvN�Lߕ�"�#>�ܥhB}K��20<����L`�r� T.�6$�}`�t�5@�Vo�S^��Q�^U��)�Z��J�]��j��u�Q3�pݑ℠4����X�^�1A@.��=B �a(��A$/Rݘ�U>>g�B墮���0�w�ɀm���u\Dh���|V��дVd�/="�d$y�2<�ܽ�H�I5[�f�=� �;�� �(ٔ�����5�����9�@�t4���s�i�(μ����,:��"Ó0z���hkul��%� �zC[����\��T��]I8�j�V���%1�J�9�����c,��*v�"��5I�k��OAJx�KzK��v��]*�o�W]vf������/;h���P	�$�m]���G��0�Ś��tgI'��C�d	8l74�͈��-����<txVeQ|]X���)T��G�"LN����C1f͈����:ܭ�-"2̯
|�
r���h��t�J1m�EZ���8�w�2���	�K�"��N��2lO�8��󐽶��/�������/}9�@N���W�y�f�}撶��s�վ�)r�rV�0��"�k�:ï�=�d�T�\��1��'���hF9��)1���I�'�MK��z����=�/>��t4����� �n�Л��;�U��/h-'��"6��3f.���{��}/�\�Y�Qc��Aħ�,��E>nE�ҹ�����(M��y�
�z%qO��F�q��mc���?�8��r��9���6�S�T̀	���pM	�4n�X�.�T9 �$5��+)���9������%��1������,0�֬�p�>ݳ>e�b�d�_�B�`�n�BE���De�~�U��)����� �.��i��B��`��&����$�F���:=�Q��4�r���d$ǎ��ܠ5u��x�#��:��cK�ʑ��䒾��a���HĐ+Y�v-,$�wwԌ�{�%O��rY�3�}[wY�A[|��$�Q�b*
���1z�P�=�6���A��6�#>�e�A� ��ծ/��Q�6#���bX%�QD�WŪ�t֝'���lS�����B21<�Ӹ�Y�tGEn��j=l���Rp�쯛٥�l����g���v�Ҩ�d&R�&o9������ڕ��_��nXe� -��D<��s�1�[K6oVB^�B��q����x��.��L�<�n
��M����q������ֲ�#������)����	����~T���m��U�yf�Z]��ݶz�P��4?��Z�V7Yo��.�9Xj_۸��_}�`Y�K쯜��Fg5�oT������S}y�ϕ�7���;lGFU�1�?�%Hp�!℀����b�OH�WtL�i�Zi����ꖇ~��r��:�]&#�)��)q��:�������Z��s��J���rq���K�{Rm�<��&Iގ��W�Q�R�)D�O�8�S�*�������f���\�.�E׸�b�Y�=��^v�AF�=��;�:~>]��˧`�v.[ڏ[��������A�
y�O�0!u4��$�r�-��ᕛ��씏
���!@~HD�㥰_���jRrSs`��s���j������1���s�>�1ɒ]���Z�T��V��Bځ����X�c��&]�+�c��}f�pT��)� �wQ]8����S����K���BP�5���&zY	�1 _��>9��NJL��j1�~�6E�����&��[�K���o�5vB�W2S��E��5���8���Z'b�� Srψ&+=�0���d�G���c�PL�,$�p�R��%�O�c���p^��j~��~Q��Ȁ�|��oI���T$��*���M����k��=,��U��T1X+rl|���Dae$A�s�2�dn�E�%�6����uT.�@S�	}��e9Ǎ�,o#l��ģc��v�z��� ��O�.��I��0G���$r���k�J�S�\C�����H�mn�߸q���WxN
��n^�z���{��x�����`V
{������'E����b�A{l�y�L=���3����t��l^�Y"d@� ��a�{��i�ʉ���%A[����RG1����
�H/�ŭ8�QZ�pN~��#M�7��H~��������݊�(��C�rH��L��O�[��r(��$�/ED�>?�Qh3_���Q���5U�~��'C~Kxu�0%�!�U+��2�����^Z~]�/ǡ.����r�W8���JK�U���l&�$�A��G�\�b����{�Yn��)�o6Ե%=0��#����l��$�W��cF�����}5BU,WX�z�b���Jh|�(:@\��C&/KN�Mr�=��,-�\�K:�VDGG�jː&z�6��V�����e��6��� �Ѱ?z	8�5�4�&�S�)	����^Oz6�A�X�k�(��T��k�`a�8"�E9��%���6K����/���y�����O�˟X52��;�@�y��,E����JY<�����;���^|��x�o��|wMu9{�W���[�ǩm��e "���Q���ق�����!L����Z|��P��*�|����D����Z��c�	H6x��$J��'G`��J)��7�I�h�7����#l�N�$�nt������OD�Q~tΞ% �wAu{E�mŜEwت8C�dDl5��/�,
X'[�E,�B�-M�F[[R'���*�*3E ��2!�����l6,2�*������������uG>��ʆ��nC�w�G9C�D�w�"NB�m%]&�a��$�q���듍���,����Yڈũ����+�Q��z�'�Az5��o+f�-�\ӅAK�������x�6��[<.�;{�.�־tsH�:*�F)c���
�����03p���������`�`M�Q�9�`��b��4�������HS�B��י�2�3��[l�kH����>M���G��O⌺Ǿu�r��Љ�k5�"�y�ۜ�@����K��X3��~��ȂU{��@
1�CN��I�pnR���7�1��ؗ� ���M�Ḣ+k�?_�.����3��*{�164�v�S*\d���}�*�n1��{�bE/Q�]����G_��d�[�B�FQ�Q�@�s8�l�A�)<�bq�׻��m��;�
)MȐh,����@���2 *.yTR��bLz��N᭘a����߆hAD���։�.��{���"�Q=����-����/��!�6U5�]�*����mt�cڣ2D�7�����4���H�c?ՒS���[�ش_q҆��;����֣���a����'����<%u�Y2����B�Q�Bwi�w�L�Ă���%�ɞY2�c,�7��~.5����F�7x36��x�I�$���7�4m�ܭQ�D??K�f,�xޅ���#%�a���GddK�EJ�	��߬��3E�z��H��A����,V-4��f7��h��8$���ط���P�?���)����A@|��J'w��aL6��\l7F����I,[Y�CoN[�5�Mǧᰍ��Ś�)*i�\�-��9n1Vje��ź!����u[i������� ]�!eK�'�6��)�'������1,�DP�6f�i����4?�eT១ 1��P%��b��HA~���*����uM�lT���j��Rڔ`��2���|�.��%P��p�.���4&�C<.<�	�;|�k���TI69� ~��܁p�(�|�ԥ�CB�Xz�b��3����'����*<E62��@�+��g�c��ς�0��E?/C��$p��C���:��=+�CĴ��#FO�G���G��ܢ8gg6��D%�d#c�;���x]�t�:���e�����q8�=)��f���@����AF� O���P�C��qj�΀9K��N��8��K{�5�OL�)6���7�E������2~�2�E�#�db�e�
H{z�-@as��ݻa,�ܔ��n����IU�D��q�N1�N����b_����O���[y0�<�AKzi��|�z6��1�����<�#-q��_�	q��z��0�I~Y1�怞�u�[���@�=/<���(y��,-x���LqЈn���iu��a�T��W�?��j��=��7&���:&h��5��۟�3b����>'������4�4&�Ӹ��qrG�Ǉ`��%��Z����P&�m�M�؏�W����<`�l�Lx��;n���'�7*E�ֶ�u�D5ۡ���f�����W���q�!�o�z߫��X&��y@oz�t7�!N�5M��O�=�s�x�C-�6V�W���ɥ~]GO �
3�dP/*{��Qb�`}�1� ��=+�M+l�����������M<pˊp�Ķ�
W ��N�iÌ��6�g0[�]�4}r7o��~�P�fv��L$zi�&�'ў	�(>F"����T�/9$H�&�O�:9�]m$�Úg�f�b��J=�8�h��EG<x�F���5ѱ&J���H��ȷ�\`�?F��)n��:+��J�3�'5S ��AD�j���+�խ�+A5D$����/Q n�o�1�O���HG��v�6�pR=C��8Z�m�����l�a!U�Ֆ�̅���.�f�;�+��@�w�1�`�Í��A��jiw���cۓVּ-=ž\����n�OM��'��AϷ��v����-^j8�J_eMZMW�WwR�W�=������'r�~�g��x7i�h�X߾H��n˲X���;=/�k�fDR?��m�?8z�нLؓAG4{�ߓ/l":�|Ǩe�:��gm?�h��D�gm���n_Q9�Ɔ��(x�zy� [����QfDU��y�ԲS���h�`@8�|�쎕�+ �Qf�͡$�ʽ9�ě�̰�[��V��9#��i�	�B��������,6n\���˅�.�֦Jx���z�5t�ƌ�
�Tq$�z�dG��
wi�װ���WS:�To�L��q3�4���o����=v�:��0n��p/s�	�[��9���7WH�"O�$��,Ï�*,J����p���~��O�_����?n�fJ0�/S:�u�k�)|q�մH能9���F�O�ډ���&��JG�%H�,|Z�`���ոN}�<�LE��Q@�+��4�@>i�-�c����?Ł�+6i{��1&�����dB�Ղw�>�.�~�H��}�}�E>�Aj�;Va֫�r�?*Z��O�g�?��<���}��d��6���7$Ns>Z�OUN)RW� b��������C�V7Hc�=�qB2s��f7��GIܳ�e�mS"�|_�]DRZ~O�wƈ(��L��H�����^��A������7�XO�d��#���8c�45L���X�z��;����}�.B�����T��]w�-��k�:GE�X�	�:���H��#��_�Š�퀆s,�P���nt�5��^�ʃZ��. _�S'����IGs���{���Kw!�r�^`e�>�U$F_���,��@kSo{�_��0�p��]��K�2EՐ5D�T�&�#3��1Q��7�/=⏛�����B��&��a9�ɯ�Js�_]0�3��fE[��a�Yy	T5ڤEFƐ*<�Z鞊#�0;��d%��Lo-��ʘ^b$�jY!}Q{��Z�I7��v�Ct�\܃�]ȓ�� �f��DG:3:�$ueـ�p�K}2�IfQ)U&bE�=b}�Gx�Sj�����
�N�)���D���_���xj����Q�Wͦr�#�*W�e�p��������a��ܱLC��_��~�Q-){�n�*o+�Zr�SZ�$�zf�� p��kբ�C'�.�u����xEB�/'Z�G��b���lB�P�F�C��	2$|���k:���D�W���.�'�e���L�7/��p��E���%�4Z4��h�j?�F(��Y� 'Pm�2��~�U"�4w8&	.Ρ���s~"ݺNޑ�6L��}���-a���\��M����u��k���j�~� B6Z�ɔcAm4�u��QOO-o���u� c����
lĈybI����\;�v�`Q�	�3�,���RG�&�D_�����G���
!��`X?���.��\��g�?�IC�5������&�,�9��V*#�����`�C b �J��-S�n|8~�����J�x_��aO�8�<�0R�zt~kЀ��JK���&�Q��S�bܨ�9g��&%&j/�O	l��W������.���#ܤS��[��tS���\jG������MR�����cj��|�'~ �ϵ�����רb��D!R��4a,_V��!�.3��a<���E묇�K��P�_RK���i�b���1����:������'* �b-9��&�"<.fS����6 ��?�/Cr�����Q�O(o�����̝,�h�hc\s�W%2���eM[kɦ�D�R�Sƣ֑�a��ձ����.��U�%s�[�%�� ��F���S���K�2 ��$��؟@�Ƨ�&W��=�C��	yjF�M������|�dpB�4n�b_�֕7�`�:J�ͷ��Ac�8#߭x�	�Ǳ;�5�jz����7:�*3�&�z G>���89�]�vHB�G�-���h��o|015>]n��\!9l���w�t�WE[	��۬(0�`�P}�F2qH�(�2�~O�6�o�frr���O�i#g�ЎR_+���o̤j,����ff���ŉ�K�LG��1�RX
�k�d���LCoB#� Y(g	��j���8�y&$���E�c��=��M�ÛcB��1�J���K2�:�0!:���V��I9��e�Y�T�co
K��I��)_Nu��}�/���:��l�p q
��^�v�P#�u2W��:�X�;�� �{8A��)Jٓd,�J�$�Ƈ@ǈ4�I�@�����?��'Z/^z��)�zQ �8E�I���	����pyĔ��5�%9,7���\�/�O�Xm��SR��4���S^:x��r�P��J����9F+�|��e������C���S�����0t�e�9=��.�Gc6o�H�&C�ގXb�L�������w��i�/����U{t@c��$vT�p����֟TV�(�B��h��8<�,)�Ք�@P�!l2g/��Z-�ԿcZ5�G���N��*)8"���r8K���}��������5�f0�5�/ܬ:�u��Y�c�d5C��FO���*d%Kg���嗬^`ոxq7��K������k���`�q&�p̥�rQբ��i�3�����F��ȠCP<�&��"6�����l|oe��`L'I�����!��o
�/RK&!"�m��/{��ʍ<'$r�Q�=�n1�`�Z�����7��v���0&P�`��*����q��-&	+;�I�w^����k溧!�����H�������K�ȓ���)Z��g�Ht�?�l���K�6L�<0�V϶x'ix$Df�7,�ZW6�.���T�z	��:�ǈ����L����?�$��8@�a�s�졌�u�k�L� `�(iܛ� ��?	�D���i�n�����cO@!@��t�AWy���h��3D�;i鰺R~�m�0�۟&�?󠄞efLm��������V)���H�t���t-`[���^Ւ�I����}T�����yu�P����rZ�kw��\H����4<�D.E�Ar�D�rQ�DN�I(�T&R�����$�"8P�n�V��n�:�iI��m��N���\����#B�4����14�e<���v�C�	9%�7� �Ra���yDIڦɼ*�u
����Ik�ZZ{�c�t�qi��nPzP��!�J<�����K�ĝI��"���,p��w�U�]|��(s����$"n�S�h��o�E$�{����&ky�4��!6n���5![>^kb�e�Ю���0��D���}���~4}�Eї��$�甯re ��3:OR�ۻI��~FT��oR���d&bX���QL��+�kW=�x��]�-��R�9�9O�׫�`��,��u��=K�z+D��Sa?��݆���?5� �6�t��j��7��J�ڥހZ���@�o�`|߰���i�| Ց橡ױӍzK�	&�Wz�qՌKۖ)'�����ޚd�j��hN8YCb4�lew9(�Ѷ5�Ct&$zIR����`�g�Jd''��>�Z�i�w�����@��G�Rx=�>u���Dw���4�#R$&Pe��Y�@O��CsO
�X�`:r�y�_���٘�q���P��EC	?`��"������m(h��
Q0�\�#��\p@!8�'<Q�(��8�.X�z�?sl�Y=�R�op���l0^~Of/H��z}�-(��v�q����cd�W��.	Ň���	+� ��4������~ �~��r���`�aظ��pF)�Y��:B]A2�o��H��3�x�e0���������p�ߋ_$�88(�j./]��1n�Q��n�����@`��2eu��@*�+e`Si!�i5LZ@R���gb�kU��߀������3(/cȀ��	����w��@�\��F�g�fc|����J�*ݬ��7���{��`nLf�.�����ż�VQ2s��yA`��:=�P�5ۡ�`���<Zi�|E�hj�����62&Ǫy�2ńϩ�RЋ�]d�٥[�҄J�LFՐ�v	؊7�����`m���֫Nk+�eR�H,I��X����2���ƪO�1�q���lq�%�
��'�m��ZR�
p���b%�%�t�ۋ�m_ �s�xkƶG��A�jKA��=1"G�\f�k�~�I���#rd�����A�=�%��Y���hBi(�M$�1<R}7��]|����ȶ��0	|9&%#��*r��m�^)���÷vPt�<���\e�45����x �.ra<�:~[�Q�I��6?�_�QaU�4=�����
�wL��G��9��*����YAS��\��
�R��3��򴪗��Ynn���J���+'HS�?�LG�1ˎ�/��2��9�}���C�"+GnAW����iH�S� j9&�2{���悏A�p��_��s%�����u������cJ�o�lp��G���Z+ܱ|���dyt���D-������f,��VD#K��I���F|�Y�$v�xMA�H�č6�,���)� �j����Ɇ����Hr�Fσ�p?/|$��v��r; *-%�X���Eb
6�;?P����
5���G~�wv?<���d��Ep�:>�����X.@���n�sS�q'Y�-(Q��~�fz_3�V�0b��O?�ۇ�b
���8-�X�N��䬬LŸw�qjiC��PƊ�rp��5��Μ�P�(�c��WϚ��.��fO"F>�T$Jƹdn|�]�3�U#Fi��?�R��oΫ�6���gan�^*��"l�u�?��V�=4S��z]�$�����"��]7��k�a\�(pB�Fn�h"7��
��r
�^��ۯ)�뭯�7�s�		~�K�Oہ��P��F�\TL�Y���k��y;��8�G���oV*٥#�ԣ����\��:dj3�;�(�z,sMmұ��E�h��b3��y4��J����&6��d]�*!�%�!�OE����؀���/��+pv��%�J+m�������кV��v��L�|���t��F�+�#	X�PBٛ��4ເ��P��w�^ꩊ"�����[�.	Z�j��b�P��@H�g����8�d�'���Օ�[�w��!o>�Y���uD����i�q����#\�$������dRzH���Nf���P�<�ř�?C��Т`u �Qi��'7�	x�U���k�ﲌ}��g�u���
�4�Ә�dܸ�\G\�� ��.]�N^��9���-�l��R��a����qyH�.�4c=@��p(2�:p�&��aY�j��/�E�;�Rx-�0���T+i��1 o�s�b0�.��I[����M�}�Obu�O����k#D�)��ߵ�]�˵8�D�r���+��R2D�T�h�VQ�^miێ��OKz�G�Am9"|���{7
�9a�W>W�ؔ[f�WӻNo%�*2ɂп�ꅈ���O"�o�ط���5��~��!d'�'���0��"��m�<�(�H��Y�%~>�w��}����y�o�<_�$P�c��s��0����M,��8&G������J����I(a�OJ-�'��K�W��MoCc���:1qj�݂�8M�Ru�� �t��)�|�2�&:�Ԫ�k�r)}/n�����/���|�.��ɏg��M%.�J*X􊖅T$�)�/��7�~�Y|��¹1�h�>+�-�U�4}Cq4���͙(��N���������P���>呖�b�1:�����OPA�R��q�'�
M����\���>�$��As��\�|�$#������&���h�	ѓo��=����@c�����_�s�����YY1������׊*��{8�h���6�ы?bD���/���d	�UuN���*t��&	�9�`yQ*6��IL:�N�̅e+W1!$��9�5A�յ+�
�0���;����*�k6a����S�Ʃ����df�ms�o�<�=�A	�w�mӕ�Ѳ>нxRmA%O�������{��9�]<�������= ���g��.��|��W��D��g��	���<g���Pu9�L(�v~"ǋ���r0����g-��K~�W�"ӥ�b�ߔ����|[X������#������[Ąi���.�|�G=:�+���?&��Hϸ���7	�^�
yGG1D���jX<?��T�Mp�+�g��i�0B�	��%⺗�P�r}Aj��p��BKYծ��f��`1�Yo~De�+�/�ጹ5Z��;|9��<`yt�-�������B���V[��wƪ��6��6����Kڗk)Bp�鯈|��Cԉ������4uI��+-u��ߟNs�ܓ.�jvH��Ι%-C�h���T׆
�XPXoM�P.1��)i��)���]3��iW���1F7��������;?��i
<��²�x#Ŏ�ӹ�5����ϥբ7���&q �L�"���w�8�B���m�P2�WЏ�ĩ�fP�	էO��Eg�Ek/�I����hd:�0�̫�Wvl�|#���Km���(J��"��b��h���`3���ů��P��2�d�T�����2�<�>�t'�M��b�c����8hQ������N�Q�������N���lHx���9�xC���z�uP7�$&�/gi�<�j��|~x�/���x2����<W����>[�0��� �}^m��pa�2��;j:��\�G8hX��$<��Y�O4D�v*ͯ6�!h̪*�0GG~H�Q��_5R�h����ss����:�6�P|^��<� ���%�f�9�,���|t���2J{�I^4x�J	Hxz
�D4���"��ʦ�)Q�LM]L�
Ο�z�u��v|�s/I���8B����	n/�)�@�gy�r��lb�:�0���W_T�W�5R���ν�7���or����"!Q��lb�B��3��/B]�I��L����חpN҄�Qe����>���O��_� "XlxVHYEB    fa00    2e90� S��y����lB��Gmi���^/�x�O�+W��.>a��#$��89�t<�>�9���]�]���u�=�#!�@��s"^V����ǻq��t��3ʫ����c����&��{P4-�/�a��>���b�v�']����f�����=���_>Wc �V�D�C�ᘎm~�����d�����8�'�8˄��7BX�#�d�t����P��|�ar^l��R�j��E%�<#󒬛��x�c�Il=�qdO�K�R."��t8�Qi�/h�O<�B�G���$cy2ztlY�\h���c�i�X[�O*V��c�ą�U&��u�B��/%�뢶�t�i uW��1APZg�J�WU�T	ǰl7�-�[�p=���\���W�l@�G��t'ظi��������W���I¬��n6x��w�Y$ŋJ�G)Lܤ���H���jҨ�o��ƙ(�uP�J�5鞱���TG|��C����J�rĎ$k�u=&z��1�E�گ���X_�UPa@��7O`���cC�9�jr��F���C�8o�e�ωT8�e@��D����b�Euha阣nz,�=�_P�����(�R�F�O�턼ڊ�(mu���X5fB���F�M%�x>M0l�Zb�[��E�-��	��+$�t�)"���4D����"�f,����f��(9&/59� d�.Q�M9��Q �O�X�jb�f�G��d�oy�u]�G �Rт"�VT������HDJ40ڦ�>"�ԝ���B�_A#��k^!�^�Ffr}��3��c�g~�F�j��(�?e@�A�
u΅�գ�t�P-W=�Tyg�װmP�ή�hZ�gL鳄�	Z������`R>�J�}���{��C���rR��95��R ���O�*&����xzپ=����m����<�R@Z��a�PLݣ2���&h|q� ����a��}��J�
&_cܜ_.1����&��<H <`' (I'W��%�ʅD1�١���Ʉx���|_��oJ|}�����!<\%�:�2� t�i!~���K�!��+�˜�w)���󲭌R��MՈ%�!u5��w�L���e��I������a���+�,����I����Gw��e{ ����x�a�h�tȂ�����Zq2+Ċ>h���V қz>"�Zna��z�S�f��=Ͱ$�z��g4����F�b���(�B��]���������zG���nZ�M�g~��Yƣ��rB����℻���}W�.��Z�ڵ8|ڸ���r������`�`���7/�k ���T����j1����H �M�j}+�A�����E�'��qG�K��g#���|^؃6�1�l-��V$z$=���;cW��>t���s��N����}y�p���AN�y�]��j)o����mT���ÇYV-?v������h{Ex��OC���tS�'��k�?�G�mر��C?�ػ�پ��6^؆�莇o�5;)nXy�/h9��'1W@���D�1�&!0T	{ I�yZ�'x�V��jڤ4c�c�ћs�Gn�|`V갣��ޡ�K�{
�7��cmӕ����;i f�%-+�cy�b���Xe��YQsT���sJ�|f;��5�f�4q�?�՜����ׄ�WY��ӱMWvR�I�R=̕�o�1։�(�*����~Ƃ�"��ܙ�� ��J��A�_��
�%�m%�O*s��tr*�Qg��'5�f�Ȭ�zN �/�}So�"�u�t�au? ���u(��K-)����H��H�]�G��w5�kk���/�q�B�;T�F�S\)^�.���7v��5�'V�Ң)g�,hT"� ��V]�Eb2�2���!<�j���
C���P�AT�{ص��k�f=_�g�|uɮ����T���|/�Qh��i��KW)^jJ�W�J�1��G��T��5�8�3�b����y���_R����"x�B�P�b�c��+��L���[�U#�!��1�6����p��Q�H��'�
1�T��<$۔�zD.��*�h"2�N�GQk!Z���Z��S4��7+�L�ޭ��Ӝ����������1-yp���.�7�N$�m��9���%2���=��*5�w��a�e�����p�U>���E:TW^F��Cj-�<�O$�z݊))���fE��Y�6�Fv�/�ѯ�D��<�o���^,��H��W�
5T��Ь~�7�d��"��͵ߛ�n4!a���*���3ٰ3�ܣ&��#ߥ0
�����k�^Lm��J�L(y�-����4K�lV��o�U�����B>��.N^�,�|��Z������:�ڟ{&�΁�S��⽲��z���e])U��s��,�|����Pw�����n�ӹ"4�v��X�v�%�o]����z�$YCW[g5�����Q�@�#�r[�d�n����V&LH��d�-� ��Oܺo\''9�P9w@�RR�c�C�ߍ�b��a��"=2�����C_/�-�#�t:��z������нb�C0��_Ԧ�����,P��H��6Q�ɟ�mƦ����d.٩�S�3��.pTSe�E���I1R�����s����+	^�]?���_`�4c�zQ*NZ����e��o�������&Q��\܋�s�C}��MV8'Ec*l�W<y!����Eu{T��t{F�>I'�R*��Ŋ���G� �Hm�3��;u��m� 8>���h��CP���A��HH��)����,ԝ�;e��rڴz�H�|zj��hº �%��tK���>����=���.�9�Y���M}*��u�;�bAm��\�4]Z ���9g/��ݲ1��*���Ҙ`��%���KV0����\��c��l�+V���
O�?���O�L�7Y�l���d��F����2둧���[���1��y�K+����2&��H�El�ed�j�J�QI�B.�w��N$ 뒹����w��H�ٖ������� �D�ŌI�t�D�΢$����^C)���I3&J=�k���8,]2|[|=,ވ��m�T�I;~-�� $[�O7Ȝxz�Ē���7����Uª���N��<�Y�5
��b�5Kw�~�"��d�Ǜd�,�e4�%hP���c��ʁ�~�#o����~7���A-�X��5����+������L����N��]?uB爎7j�=��J��F���2���Hp�;�+|�c�=[��E@�~v0��(�^XH�1�3�a�s��U��,K�霉2�~�s��~��$�!���ćhMI�+|n�/�"o�ǸHWK��ۀ��SL!�.}Ň�)�g�Z~��̺���gY>?&�X#6�]Qfj�aV�V�����|[��yЃ-�������{�d�/\�B��\�Q��R�(�bI5ހ�����p�E7$L���[�v����y>]��D�*�����E[��1+F0�e�0�EľXp��V~d������i�Z�8Zx�T�^ݧF�K�Vƻ ��~� ~���(�Ί��=��8|��~������8���n��{���Ĥ��\�.��-�dߴz��ӳqKk�?9�L�Ɯ0�5 ,;�r�煠e��%���h�L�|�m��@��N�D��l`�υۇ����%�x�6������qLF0��5R�^7���閯�h*x�zS[��yi?Y�`��{�	���采�X��	�B������:��-=܉d4�R,�����.�UG�^�U��d|�0��E>�Ɨ9���(8N�
�����Qw,3�����#�=܋X������Q����w�$t��S�ts��v1K4���m(T�b0#�������Q�Ӹ�$)�Hh�EiE��C<⯞�B�̱k1����3���oF|��=&����M�ݪ~"n���"ƶ�.Ƨ+��穰ҏ��?X<uB�)\����:�L��31�P�o�j2͖,�M۾�0�z���N�|D���q���F�c��{#)�/k���3���"�ǿ?��RDp�\�(S(/u�:�
.�~��s�QT~M�O7)�u���1'�r�"�kH�Rn�p��}���̺���B����k��A����`�v c���5��k0�'�e�o�W�ߛX��^�P
	%�%!۝`��Ǝ�z6�k����bD{�-bf�/i�P������gU:Y���������E����b��\k�zϽ�9_4�M�>�H�����D�%�N� ����ȓ�.ϭ���oEͱ7��ѽ�m�>��}���<ɥ���o�k�Mn�2&��V��}�,�r�����-�9M�	v�Q���y�A*�ĸ�I;�m�٦j�`�2�SX����\�	kc���D�h����Jz�ox�K�r���
��n����įk� � Oe�$�
U�c��8��:#��Ċ�`���[n�����C�*��z�E�U�&3��	Tx8���p,���U�d0B�Xr���e$n�Z��r�4ˌ� ����<F
�lKY]����<�c���in�l�co�ju��c䡹�f�j;�0b��#ĭ׭��#AXM�[υ:ݟ��D����݄�~mNeQ� ���1%Q]�V�Ũ_2�#�-��I~�N�Yl$W���؝�[��s~�$��iҎf��Kt�B�Yy"T��.Q��1P�r��`��8Q�T%��{G�!2zm�*��dIVá���z���TN�GRr�7��Ѩ�������DzU�A	Nꐟ"~�7�;p����a0�qh�%�q3v�>ɇ2�����Ӧ���*?z�U�v���Q��>��'�������[^W��b�c����JO72gp��� s���AQ�\J�w��Y�_�c�RP���C0��9��'z ���n�g�t�-]]pP��
1�_�V�~���%Gy�
=�Bكh���,���θ�G����r<|�?���h�Tv�s�ɗ�(�������?�����N����(㜜��-�k8�Zb���A�:r��&���Ph*�!�}������G��2���w&-��)l�0H;�i͡&I�����R�����QY��sh@�)��Yp�_�H�L��#��_�������Q����{[�[�B�Sj�Ǝ�3?��|��u*Zľ�:��y��
]2����X��<(x�$���>Y�0�[I���8C�/��}	O��Ǯ�����hЙ�>E��Z=��#T蜙bA��r>SD�ѯ�b��$Z����v(z{�2T�y\x�����U��>�}���@i�D��%��)�-�x�����$U�y�*�4�P�}�/R{���u�ǀ*�p�éC[��48=��E��7�V8A��h"a�⪐��@��&������"���:��f!#O�H�7L._㵵f	Z�>�)��9�
J�*��_aP��Qo4������T���� t��m����L=1 �����|����H��=���ASɑ��:�|�-w+�����P7G4ig�<f�g<�0e��[u�F��(�Z�u��'��N\<��9�q.4RO�!fl��
�����E-�	Q;��Ȏ$ӓ�_�ȶ�3�%��/;!��^+����ո�ƅ'i?f�Ll�ߓ�JYx9� G]]�N��WZ��w��XF�e^���+�X�&w���3�x�z2z"��{\C����������,r@���(�E?�;V������^���%ꍏdW8_�+չ��e����
FU�����T����e�W0�������#P��|��4*I�۹	=P�����:���l�����#�G��M�4'������9<.!�n�qx�ZQ[����4�4Wt)ڧ�X���v?�
Gg�6ߐ8��`+h�VR�ʞ��F8�=V��Ms���v�CzQ�ы9W�_�~w���k��?��MAe�#�$�8܉<�O=q��o>��d9��@�Cfᐇ	�	}����&���r��ffZ��`��@�P&Z�r'w�:��U�!s ���V��-�%g3Z��-��x�����$�|��ß)�����5���V8&a>�|C�2 ~-�@�-ag�c�n��@��L?��a�@�˕�^���]�ܵ�s�u��*q�#͘}V$�Є�m�3
�T�YN�&|��j�a�]`~�A���h���q��=�=�x`���V�za�U�TdM�cu�2W�V z��#�ʁ@m�3���:�`R���A���ϣ2��8��D��yR�����X�̾�)��~	#��FM@��i�p�Tx��V�័Y���sh�̃[��OSQR5�O>���:�h<dΰ{�q��Ϋ&��r;M���0���~�pFr{�X�V}R��bq�hYӆ�����uFEw�Z��h�/v��UQ�g��1`PM˛��&M��cF��j|�[���v2�bG�Ȼ��KP �N���]�j�};�n���M?M1���ҳ�B��;������U�}ΰ'>�Wu�������3�;~'�hUAX����T����"1~@J�`hZ��={:����.�e�/�Lצ��x����1�ky�r�ݮ�aT�^�cQ݈4m������������H��f�.�켅/�))t7i�D��(�@�Z2��U��v:��K��^��n�
�&!k�G#��?YWj
��)�����d3�~�?��7���:Jeg��P ��?�i�ȾH-�-�D= :�;�Ѹڙ��&��?ćH�F�R��$g;6�����rD�`���zeO�����w(�>3gWL� g�����܈����댶���lIˊr"�ʐ�����+q@��o��_w �
�'9�'�.Mh����Hbu�^��@c��|e�HH��ӄ�L�'���3	��թ\�Ϩ�pf��ڻ,��� �E�������X��ʛ͒&���*��h�}�b�[J�(Us��A�H�LN�|,��A�69��/M(W_U�L��@~��8��ԏ9B�$qu�&CȷYgIy��;MX`������q����)�e��o��P�]�jW�Ҧ�R�[����;���)����:�)�\���#�A��%����o��h�h� I�B��b���ѢѓQ�u��=���^}oK��=_խ���Q�E�#y?�Gi�d������҉�M,�@k]�	,ү�{g��#5�C/��}鐇��\.�!�ɀr���Q���x�-1�%�u�"�E��

���Z�"w��I3���ei���]S�O���B�A��|ǖ_�Fۋ}(���8�ߘ�+' G�$�5���[�pr�h�������0�� ,��Y��	͘�J��`hg۽�X�Ҋ���}�H	�]��u�:����t#Ύ���/۟�׷��	���r�o�'���{(~�#�M�(�h#^VƳ��"���oh��1�c�s�+�M���5-+4�����pE^�d�,ga�@�7���^NQ|�8��~�`k?nb�����fwW\Hkn�+&v�;}JUj�L�R���|�~���߭U�ƤֲE.*���Zq�E(�9|��<��]�]��x0Y��h��Y�p��J��;U��+�:�Y|����j_���bk��!]?+�43O0�9�7d;�H�y#hiz;L̛����\�6�(M8�fF�|����HD>�_���#��bS�:_!޷���Y�?��q�M'+�8�"cM�O+��8��X�R�}���v�u ��,#��y��ϼ����;#`
l�B�α;~����S�Pέx+@�MT���z��;^��&�⢏���LQ��.�m�����%�'�`p����U���a�0�)�	�V���	;A�f�̰0�F��gTd�.�,R��T�a)*
O=J!^́M�"M��Z�(����N����#�$�^���B�]�S�X�y�N�x���+���2��� �lf�sb��{��dQ�O�|�"�ӌ����N@�/�oa�Rw$�ؽ��`�,)�����/��ӂI�&vcҾ��b���(����c� ��Mb0�3�4�D�CL����t1ә{�����l�3�\��k�t�r�R��ي��&y5%\��z�Ǒi���fI�67�P�$��k�������E��X�����@ձ�+Jt��X��q��Z�Y1�+�h�a�Fj��뭧���_}�#oH����r����'�TK����z�G�"��ͩ�Y���ݎ�5|�?!�𧚃/y�v^�l��"�Mu�W�$r[���?o�*m��_wu!��{ NƠ�C)�`�D��ř��[��V�b��Va���[8���2i�xe�aH�x;�Dfʧ�2^�DwJdõ7�'��՟��wI��^����6��#��X���i�������m�Jlk�u!�g;L	�`HCy�z�4N��I���
�$���п��ʈ2�^q���c�O��?�-y�S�Mvk{�F/�J��H���\?X�B}�=3�/fP���z�?C���H�����sxI'ٳn�ޘ�J�Jڂ,�9���P���� k��4�e�_�q�3��4J_Yx�HTu3��ߧB�}��%�1�a�,��8;J(�Ô�㡥Op�ף�,i�!į> ���+a͙����uX�������f�A��B��f����2�5��Uo�k��,M���cz��0���p�qҖ��k�oI�@�KfV�m�
:��3х>� 49��Ot�ӾH���e�R�c�������Ad���(	�^�e,�V?��v����d0������x�r�p��\���'�f�����/���X�-k���_46��,roWg'��)��Z`wA0ȕ��b�)��_ۇ��Ȟ�1�t�[��N-���z{��L&$��R�P���������i�u�(�[�����<~Q㧂Y1�sA�[I��[H��΂�Ə���-B���}��&Ը�B@:�
lǛ��9�D}	F�#Ⲋ�v8e�p �2�d쿄Ļ��
U'`��f�`�qՕK?�)�a	Dy�gNrF1�6� ���ӫ&^���6�á�B>g�n¥�{�p�lgc��t{(a���ݧ�@WޮX�=1z~V$���
J��q�4j��;d9��,��0t��Gl�@S�|�?j�\(��k�Q�;\H��A� P���,lA��bJ�)�ֹ�պ[@c{x*W!�J#=r�J�?_�D���ۿS�~ f��D���8��/y|���j��0��
��A�� onI�<��t����r�.�X�j%1�s��J���]�Τ�[>9���QĆjM#&���ɧE�4'�7��Yr*h�b1�Q�Y��=��?)͔�)���s_G�;�������/:��@%�r'a�~[E�S��u�IR�췋��x���mUA�]$�F�
��Sꢧ��Ƨ/JE���=��y>����k{f���&$�,�kv�u��_)C��ώ��6�ǭ�%��o�%��7{���6-�-����R��R����5WU�'�L�)�#+\E>�>X�[m����,�؍0���M�S�"P�}�po&L7�r�s�B�[����,¹�mJ�F�K�ƛ���l�|
n[�l��os	���:��Uh��H$��S{hԼ0�m;��}���v�F��-h�z_��u���%�x���;�z�jP��@cx�{Ҫ麢Q`�/���b}�-s�D�p� '�x���(����eQk֫����7pU}E�'�=gԬ��d~��u�'A�w"����Hy.y�����O����B����Fa��.����w��&���R��f�M�L0Ì�-��㓮�L�X��֨��-��d�P�T���O���{��X�v����v�>��n��߽'�E	V�Ύ��C���I{x%�7prm1#P��\�a�kN�[�x��暈`��J�U�-�M[����Tf�s A�o��Ub҈��6} ���n�
����mH�i�Ys�+0��*@j.�a����6�l$<�-\pЃ���)� ��N��KN�h����(����g*(n��$u���n�a��̘�{�s�n�=g��N�@��\�ʅ��ˡf��CtOX��`��i�ʠp�ȍ�@䧌�������2�n�U�<�_ޜ:��;�CZ�Q�c��a�%�͵�*���l+x:"���Cf�V�t��S+�T��Oܬ` a�	�%>�	AK2N� y8�>D4)�ae���C%�Qnk��n#_��P��"e�[�C�^>x�Eܒ��I�����V��Y�T��EGdv��}�YH������Cb��B0X��M�BĬ�����ѷ!��z(D8�:��U$�����d&D�i ��ci`Ѕ�ՆC�B�y�C���o~&�H;d'%�H�!�ڨ�n����X���!�o��  l�g+��\�T��#8�.F!�������z���#�#l((����󽬗���P �l�2`��Y�BHCŒ�������d�(j/��ۗ Z6}�]LN X�ۺ����Bwm�xk#��s����ᤏb~p\�/�î�(�|6���%�c�F��i�C [��=�; }1:�R�~]��|�w��N�Ԟ�]����*�Þ��R��/�zU=����c���yyҗ9��#��O�ϕj>8��Und���?��vɹ���;�M���H ������t�x4������㟊ִe 9O8�e�/-��6�X&��듙$.?&���#���|��=��|����iϲ�(�x:� ��F���l�@^� �*�#��e
"�qlo��S�VUt�vS\M��{�'Ꭻ��n*�\]R�V ]�>Z�k�@�@�i�P�kT�����"���"�}k1$������7dP,.�� ��	o�����/��T Ƽө�6&Xp\�Td��Յ�O���~MP�]2����*M�������E����Ѱ)Y��Zf2�i�!n)�j���;E�oK�>Rh�w}0������%�k���sgv2� �vY��t�(���Z亦��q��%y���*f�p�� ]��_�2,����k����7��78��)�#�z^�G��*�o&�8�@\>+��]��)�%�7Q��ab
(C+z����O)Li8�]/�^�ڒ�
"�9�6�ݎι�a���ܥ�p�B_2��
�z�]�������E�]��y�&~����[y}¸6��0��H����eR�7��m��w�&��y����g�cʒ$�;U�]W3��	H�����FJ!�2��̘���^�:U��R�����N�1�5�.�{�u8���	B��HW�p���e6Sv��yY?4�:n5|MT�A�?��͇��^� t�iI�A�}r�w3�`4�yF�ǹ�C j�2��항�r�j�vr���¸�g�<Q���v5%ጂ���cH��^^T@P�����̣ !�u�h��z�N#�l�Lb$M8x.kȝ����EP��V�2ci��U� |�k��U���r��ך��:�T�eE�5F�s���d�j����*�^�kO����*U���qX8���c���1��)	p��y�_� �X|_��հq����r\����>���Q3����:V+�`A�dG�ȣ(�c�,�2�W����V�yc�EE�4���I�Nj�I-\���+��,���F���Q�U[�)���fyw�Y�rp���0
<�U�o�Sdy�"x{�7�kt��uP:t����1wS~b�(�s?���+̔���}QA;ے�4t����u�J�I�C5������1 �� Ů������75�\��S�CF#���~	5K,کN�[L�Q�w� D~]WL������P���i =XlxVHYEB    9e01    1c008u�U_��[�G�ѻ��%�;�
�1H,zY�f�*k��ǘ��s��<�hw�Ax�2-1��[�Q�X�?ʓT�|���^	t"�!#[�%��-��898�ed�U�U�� 1�Tӻ�o'jwg`��'��7ˉ�p��G���rw*��y��Q��]�����A�n?IOM��J��^|�$����ʫ�V��ߑ��0�A�3�i����9����iP#��=��aZ��9|��aA��� 9~�-S��xH���+�b�C�mR��i}�y���i��{X(�I��K��@0�ᯃ�����J�Gf�.��~� 5 `�-�K~
�2zgI��Iy�Em�/��+jn�e�e�������׷�"qlgp���roc�Fj�p"�
�Y����an����|��[�	�y�jO J�=w�;Ov��xa�<[XL�o����f ��~��k"o�w���K1��������$#�ge��$������6_�V�vt?��]�CROf(����aL��*���|®S��̹n��iO<���;���{���(�!��3_��AT�ih���*;��=�h�ቓ���z�U�UҞ� �/W��x��=��)vows�5��	���iywG��Ncu����^�n.ܷ{۵�Q��'�Ū 7^b��N����IDm>�nZS��ql�n]H��w�~��MJJ��ǥV<��!���䐣0���i��<�'7�=+�9�x�~p^ �s`(C��Ҹ�H��Lv�[�	>��l``�ܸ0��H��ڕ��=��L܆��1��O�+�8�1��^3C�$?�=���>��:��U�D�A��!6��a ,Ci�N&�0b��_$Ǌ���@����M37	�M���@�AT�l�ɳ��S/\�/8J�|Y�S!.YQ>�`��"�רx]�"P�Qq����C���:]di����O��LM����꾂ҽY?���c�1�ث��[�58D������u�OZS1��9~��ޥ:y�w��Ө���<ED�G�k���Ă��J�~[2f� ��X��a@�bx������I_eI,�޳��8���K	�a��?��)�`�ʿ,^�wR�z�z*��O0�b���{u�*=�2.$	F�NX�,M��>7�Nlg�H�O#u�GI7v�w����D.Ƈr(k���ͮ��3/:EEC��xB9'<;��3��G;��f�x��i�j�]VF���2�̓oYU �C�bTı���߭��C|�|b	!:�h�H3�ZǒOe�;Z�X`9�?��1Dֵ�%д�S�\�^(S����-�m�X鹚�j0:ŦͱD���~�i�&#V�c�W\%��81��LoA}��*�"���y��:FR1�vgT�f��G�#�3M��J�FӍ�+�U|�v�k��C<��p*Rg���H�-��6Y��(�C;45�c�;�g|A>?�D:�#L�, E+�t6��"vg������4)%���QiD�\HIHJ������:�4$�8�u��!�$V����5����&���Զ�T�l��n�>s�-L�U�l0b��sQ����+噶��F��`U�X�L&`:B�M�N�u>����MM=(}�!����sH׮�d:w�>[��
1ZF;�K��+�`b���a����i�^6*�V:�9NRh�&H�U�����������O1�%��vA�Z��nJVьL�j���|G� 8�cP�	�d8�e�R��|�Z� Z��|$3E�=䟾(w�)�GPz�8 fyA�Q1v��ȴ�Y���r���W~\���������ur����uen��lӢ�d¬�7�`l��䐻��27�mm@S�5}��5*/A�.�� >s�s����?�.����vm�@��i$�e�3�à�����*8}�i�p��[R��^~Hݵ
��&#/ �V����E�{��9`~�GM�6��t9�Cî�BICh�[يm7{�h��i�5̷!Xjh�U[�T�Ʋ�v�Ŗ�=+�^��q�u�C�S?R5��ڸJx��-��hf��wA�2��gF�O@�>Af��q�GV1�
e�I�P���d��(uP.B��/��Yf�=�,��@^�Nv#��G��{��ҵ�8���\ͨihyXF�N.$�ӎ�$i�F�5��F\#iѽ_B9�fD!`iʧk]+�����*�V#�ZI� [^?%x�F(�"A���<�K��1G'��.���7W��Xv#�H��D��w1�ʛ����WV��s��+.�qu�|H�������P=���S��u�V�)c��p��xoa�f*|(����g���s��&R��J�S�0���
�	`l/6ꃓ��Љ��Δ\��%<��9���O�:�BA�pUL9��ĕ��,#��u�^��]n�S��} ��;z���J�Bn>hO��x\�z("S�'3� �^K7m�qƹ�+x��܂��9} 9���ܸ�]�G�f�#���KF������[
UmP�cH��5���"�kDr���⢀/l=�I3�kPMe�<Eo^9��+30��S9=��]�Q���֡g�bM����3�=S��m1]�
�W��ֳ�u��$"�Xp(y�M&��l0��L3%��B��3���rR&[��ƅ�Qnvw�>7�$��<�?\1O5�z��>h��U6e�d�AY,�IX�eZV���/�}E��H��nۥ�d��ŝ��{���g��L���O_e�mM�8x~����0^L��>mv�tE0I�:f�<��]�َ�

R�rc\���c
w���_@���N�w���3F8(�;`����+˫��?��׶9hR�f*�E���bT �6�.�:H�(A^0�<dъ}+�x��Yt>���0(c� Y�=#
% ����d��� ��G1 ����*�!�S0$�5eF�{� �� ��>d��s��<����VM��f�4EI2	�DO��=
����r�y ��y5�*y,����tp���<"�U���Yn1 E+�RC���ë���n �� �Fw(�6hʏ���yVPS�e��J+�*������w��+k�_�e德^ ��e���<zG�����{?�5��p�?�$���89]l�/�I�}?�*���H-�O;�59%hڛ^Z/}�
{u(�w�jс�|�D�}����]���@�u4U8���F/��Td�����֚���\Bv"k�}U��}��^���K�\�uz���iY��a��j)Lʐ����u�4Hv$�������c��EE��(1O�B�\����#қ P�����OC��C���]�6�A]���)��n8��.�?ޑ�D��#fZ���mDͼ��e��,s"?\QђnY;��r:��:qH�;�)�ծt��mt�G�<�?�ߜ�t������(�=���*�%����ݑ@�&a��O硙 �P�j~�W /��3U&劉\�9��w��x����&v�-�� {��9U�)_��=3-���bH���ْ���'�ZO��/�Se���� o�@�Q���]�g��rOAA�S\�3T%�p��`��B��7�F���䖒��}��p��:������/(�Ky�����{a�0��]�;�FA�Ӑ.)�Xv/S��
�����_�2��P�!l�_Buñ��0��9��]e\8m���X�_���iJ9*pe��|��Y�?!A���T���5{(��e�NI��r�)r�ٕ��le�6b,J�|7A(�Q�΃+�1��s�%q�,(*/��OP1�/�!{ o}���x��3�ò�:h٭���aQ*v ?f�b�~�;��I?#g{��6�G��	���
*�s���<������B�z�1��ވ�-{v��)G�A�t�qw���m9�^�O.��#�c�i�&��q�WџbLh�2���R�8�`�z�a�*Hl�t<:��$�@γ�bT��ʹw�,!�y, ɺ�T�@�#kC�EԬAh[ݟN�T�J%���)� T�F���~kP�b��ɛ�aok~"8�uUM�pS�w�A���Q����U-��^UU�q7P����x;�%i��Q'��C���h�H�o1@��cj��yj�˦�g�&��f�����>����%���C�U�Q�-Az�����g��!r�9��=��	�ޮ�/G����]9}��Pp�AS��>n��o!��p�y�� M3D߹�$)��5X\7���	P+��ܤ��u���v�w��C�����X졷u��.�=zm3;y�Eu��̎�)�w�y�G�_��=�$��uw
ΐ�?o�.ESg�-�/��@/���>֘�Ir��?bM�r]3%C����ä��z����AҀ<qD���,flV���e_Ik��Q)��E�;�;�䡺���-[��'�/��+w3��`�ѻ=��Pc{A�h���q��|T��\�G�{���(mGRT����j��kIs鉠���O�`����������U�,N�nX)�I3�(��G��j����֌�ģR�R�Q;a�x�_�K�-��'�A�.`�����N���z�Hܨ�;�!g���	�ČE*{���oBK�g兤�]��u���oa������2f����~��Ӆ�������p����� �1��܎�A=%�k�����t|��D7�$'ب�� ���f��;~��eq�l�W��;�}�6�[}e�G�Q���y��5�r�� V=m6���x�ݻ/}�2V=��m�	q�]ݫ�L��a|k��<d'ZP&�la�|�i5���}�r�����b�w�˒�%-���=�eX�U�̋�J��Z{������F_I�u�WP:�t��T����z�H� ;�&�!�lK-E{,!�Q�צ�����MI7��|6jY���%�R�	�3��fy6)��f�ʍ�#oa�7�l1�<����OHh�qX�t*�tr�s�&D4.NXIx����@8�*�&�X�q�7���=Q����buj�x��1��.��ަQ���z�׋��3Ck���{��ȽBu��϶��i!�.TP�
Y�٬ȝ�Z����շZ����BZ�Z����8�?�ڐ<rbx�����j��9��uΊ\�780@�[!��c��xA�[w�~8�k�ޛ�P�<�Wc_�B�f�	k7�{�B�>$���S�q�����4�������;�����F�}b&x�*���;�7HO����:�%P�o8l`�<Z�� TUn�i45��`����-��,/Nq�YRk3�����N��U~Tl1��y�Y]�e�߈&+f���/M��zԂ§��% <���Y5��?����G� m� Oy{u�W��
c�}'�Zo�9��:|����ס�
�_,\�0���$	�2�&=��&kO��� ʹ�9_���w�e0E:4G|�R�e�7�u�à�sQ���x����t���QE������|A�%���_���C%���1ґ���A�wBF�|)^6M^�ɱ_�)�O�.m6�(v̷����t��88��� ��-��W;�Kؾ����ԛِId(�ϣ~}�y~|9T��tb��AqC�cWឮ�N�~1����4����+EtH���
�T��̎z�d���u��d���)_��������m֚�c!�@�3b�������;ʝ���!��d�DLPK���;���)�:S�x�]��
Ǣ�T�od(�1��B5+�ؠ��>}���}�[��],��n6�܂/m^>d�*�W��[���8�۽=cyݞϐ�&-|�L7�.��]�ǈ-���'G�D��zX�;�F��e��w��M��\�����j���85�3~�R8��g���l�B5�'%/�(�s�o�		R�����W'e���WZ��t�]*%��jEh��l�?Q���f�r(�E���F�� nLju�����T��<Bע�;���U�M�R���w0&,T��#Du7��&0��7с�A灵�L�7�����`��c�m���Kvp�nc����>�A|��y� D;<ɓ�˲��o��*��@��{��}��3����x�:�U�c��U��4�����6J�5�&~�JQ8��@&���"��״�/�o���l���W����>�FG}��!Ƀ�J�h2�y�b�9Џ-���Q��4jmƟ�:I���=)�GW$���IN�>�ԛ�T��"��M�ir��B��-��8&�s��d�Y ���²�Q*`d��H��`�:S'�e@�*OwZh��OVb5ju�����BW���J�`��e�_��=�~f�d���q�e���i�du	�:�&�s���K|
} 8�#�џZ;-bx�`:қ�_+خ���z���+�����wIA�(�)�Y�Ͱ✩�U�H"��͗�_j�c�"�ԥ�\�jI9�>��*�`
�,o�~�L���}�Y=D]�p#�����$"��@#K�~����2�Dߦ���ȗ5%n
d��Bׯ�l��1��B�Bҡ�a`q�����ݾ���Z�|�����y��=�4y+��P1.Y._�)�id6G=�`t&C���W�?����~��:~�U}	��������>'/�����m�u<Q�={�8|��>�d����A��aBG�I�&m�{�`��+�x�?�0[;���˭|�gNO�
���eb0;pNβ~w:��Ж?�VP[6nRzn�O�2}1����,mjEj[��k!��8\���\4x�$�3s��G�.@�aueVq�J�C�� �����-���9?�ʒ� �ɡ��E���R�e(����l(����EWp��u%Xk(K���2G*�otǐL��y�%	�6JiP�����5NC�[��'��~�>��,�Z��:{��Q	#9�ۊ��=����7/D[x���ig% �饽��-���*���y@x��pEyR�	��DW���q�NJ���q����^Ө2�u���D'vB%�RM�\� :ZNt�$�%+X�.����z�nB��#�FyP\����`�I��b�3���`��+�#�,u����&�1�G��T<�a�u����k8�t��ŕ�;��'>
�����q�=RE��d���dY�R�O���qG�q����H�h$e