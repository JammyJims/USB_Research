XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ���E�E�I��W���E��7WcM�T�#����(�L�Y'���DC��+!���P@�S�+a�N㶴SK\KO��t����c�y�(:"�yQunW��ׁ�v��K��W��]���
n%EøWG��-\�r湸x��z�L��'�(���C�6���;R"}�N���h��^��KI���T( )_� K���\3������9\��[�ڢ������y֍2p�!�3�Cc�p0����뿥�.��؝���B]�c�{�>��X/�_���K��J�3���**���<�g_��w���:c�c)-�-
o�	CW��hk�)\�G c�Ό0��`P�_l�G�&$s�YP�u���oU�O�I���(J�����ē ���M8m�	}G���� 0H.%yS6")E�S���2E����I�G_�����>~����u=TM��u �!`oF�#�����@oT%�������ُ�2��\�����`�D��Dg�r��Tϳ��eJρ	Ǫ6��4��"�s�F��?y�������49Jf~��z�h(Ä���{���m��+��%t[�ϙT�A���u�7:<;�g.?����ݓD"I"
Bߵ�{��W�{F�	�KK�. ��.ٚƦՇ��:��m��Wߵ�;H�6����&暥0��)��1�PH*N^e�wҽV�dv����qn"`��Q~K��.��)�-i���Z�;Sq�D��6�e��x�WfS
�K3¡Ҍ�Jɺ?[��{�����P�U~XlxVHYEB    4345     d30k=�ja�<GΞ0��RxS��- ��:(t$���|F�r�kɤL1��e����ܴ]�TH�>�0��[y�`SӇ�d\
��l{D�G�)	�VlN�% R�1k�z"qֶ4��[E-j������fJ���A��"zH���d���꺡�Hν�&��7i��Xw�[),��>iN�"60�a��\T5��8\�ob���r4$Q����3��!�f�!qM���z��'�fGX:} y��:, ��pqYC��\}V�ňU�bѳ�����BP���d��m������@��$����}�=|l���0j��r�M�׮��t�3�ٍѪ�����l�dP^'���� N���,X�%x0��h��恅D%R���,/�����Y5�}�ŵ���2W��N��6"�����%�1���)��ΒEjL�]_�*E��R]�AU�V��L������g��g��\As��O�XH_�j�'L��r��j��P��l �G��9^ňRKRˊG`';��޶4B��ؓ��R�����/���Ak��!;x�\�W�L�+���*�tM-*Y����ְ�Dkpׇ;�8�Ƌ<Ka����vg�j�2rO�~�i嚸�f�Y�C=S������n2O��
��ׂa�8���!k��zi9�9:J*	��}ݼ'���8�+�cN�6���5>���i�moM��/�'7D�|uA��/@���}yd��&���j>� �"OB�s�[��Ԭو�Wx�)��[����_��}��}y
'��F�ǽ�n0�o~�F�3��WY��F��)b�Ȉ��zc����3z�����=�'Ux��ӽ	��5���~Ӛ�}Pa��!��[@I���9���/�axF��L����Jѱ�b��O����r|w����=�U��)�a��Ξ_z�%У�e2�_�s�č��-�����rj��:wMܦ���gZ믵�&��[����\��i^�{����u�,�eg��Ta��+���3��b��ˍÌ�H!�>[��*�S{2�M�}��Қily��r(�ϓ?�b�mUz���n�}jl��!>BtП�i����|�BWEBf����p+@elp�I�� N6���Ry�	9V-����SP������zj"b�
9��\��-��!�=4�B�<�G �5ⓒM@���7-�+0jq��;�*|��T%	�2T��P
U�?N���(�^c6`�"÷>U`�����+[�K�3@�2X��+�	�؏�n�+�*D�dk��^}"����my�ѵ����!	:3Q+�#�m��?`(�#�\�c��[��OK�)"Z�U9=aDr�xZ8�p�}��×/���9���0��Tȵ�[N���gե�aN�q�Δ�c��w�/׶=h��7�UR|��\�#)A��s����0���ő���Ͼ����b��3�K���pf��D�9M��#2B���x����0��'~�oM�ݧ?X�HVI�W�=���;�������A��t��;�����)��Ѽ4�i�g��EX��Q*\>\�u�y��3�ga�T�G��/�
�Հs�[��֮�L�z���{�����5|r	+qqe��U���wi��U��1�͈�nK�M+�py��9�^����vzRx��)��D��[|���n�t|�k���e���j��b�CbGyߓ3����㪫�45���aGUP3��L�H���wwģ��ug��Y.�srv-(r���ǂ�-�=�� �/3��* [7s��4e �=�+�D+9��g�]PL!T�j��"�w���{�#�E�s�� 8ٹ��y�@�@�&�^֜�g�H�������}�ĵ �p�&<c�S��5�Ъ���e\P�S�Vgi��x.�^յ��Q�0��o��Hk��m k���4�����3Rw'f�?���=��"�\�%w��vTg�-&J,l��;��@�|��
v�Y}<�&qk��̤�G��S�'�=\ b����[9R �ԩy�u�:Y�žI���4�+W���)���;>��p5��Wx�����3 20+h�c�2����7tuRL5M� �Od����Q���Kѓ?��z��a�0�`�x&�P~��Ի��8���76�$��q-W�����(o�ԀD5Y[�U�%hN�-�t���M�襳u�]����,��v%��>��VZ�|k� (q{�g�<A�2�6bV�/��
��i�8Oz�&ǀ�QT����#�J�,m�,ߣ6���������a8CW�W��7W~:���)zE�7����<&i�* � C���X;�T2�GV��5N�6)��
lB`z��N�����\�ؗ z�<����?�j����t�Й��,��[`V�H	@�k�:T�����- ��j�}C�!5�����Xn�q ��y���ƻ�T��d$Q2��&D��ߚ[K��\#�^�2s���s
�r�]%��x����,����Vi�g�vN�Dfz�`T��/=ww���?��3����:/��Ԝ8���y>��O�ϧ[���v'�nTjO5�=6 %_�
�mV��77�����Z���'�!�9�K�!և{K_B�(�YHx�� ]_��੖�
����'��	����޺�vb'f ��e����Q�bWc�y����DXb���3�Q�[D���[3x���i��`�o8��4�-�K�o�Q�z��+r�ȿ8L�T[mg�E�3��J���й�����y�;6Y��Ӄ�!���K�����d@��Ex��$��G%���d]���Fu�˛J���<O)�4��$���wky���!8d!�bx���k++��U���Z�!���d��<z�V��<L� f)��ߝQ��!�P�X�����p�eg���>�W�{ 
�ms��il0���	�Ps�"�<�Y3㴻�²l�!O9 �1��U��x�K�XP�QI/c�O4��XB����e3,Bff��;Q�����K6�M8��X�?��L��@
����FB���Qz<��e��֮5�����J�ʻh��wB�q���|!wָ�ܪ��Z��?��!t��
����iw���.T���$9(F	fI�FCM:��:��;�� j�;�S�����Y�2����A������� ֵJ�� �($�K�T�{^2�zz�`b���z�3�@��:��e[����,��d3���U���fKv��Ã��򙥥��A�	���2:ƹݨ� yC�8C�.�E���r����5_3�����q똇�M<W�31a�=-�Y�{��s�^�"e�#�i��<#�:�φu��J�f����