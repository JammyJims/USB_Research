XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X��p���,�D�B+�$��)qޚ�\X;�J��z,��wұđF���ٿ�~D-�/f��>G[�r?�y�R��T����5�T��~Ɏ�� U4k����䃽x]HT�-4_��&��q-v��*��j��k�t	g�o��������?a3��~	.5��d�aU�@����[8o4����n�"G�.�pRo!��ȽQ�a�I<�7��.ʐ�'��8�;�w�B��aR��E�r�LP@�m���e��hk3AZ�BJ���Qxr���z�c���؇]�$����M��.&I�%H #ul�V\f�����Ӣ}�IX�؝JcႦ���׻�]#2-�=��|& ��)�Q�{l���I�2hS��}�%;���t���b#�ԭ�	��d�5^�����&ߋ�$�����Ua�+�H�*�D�e\�p)�.����ʘ��̰������$yH�Zf�&��gVW[���J0Ֆ,�����,Jq���7�ԋ��Q�`xƧ��Qł&�դ�m�ʅ�[jUF`1�{�i�C;��^e�hp������Ę$���?���k��h:{��5����t��O� n�%���J�5՘���J.v��NJ~d�_%^��-c*�dG�׿|F�rʄR�v����J �������;�YR_�{yp�ԑ��Za��A��&��Kx<�b���y�CU2L�����b"��YX����N��n`�O������Ż�?к�����	����"�[;�Vޜ��Ҿ��ƵXlxVHYEB    545d    17b0Ǜ�;U��H"�@��3��1I\�� ��
��w��=�����@|J+��7(4���������?�������������L'�		e����.ؕ����w[ԶF`o`�	��_��lP<�y.=c2:B𹣴�
��N�mK����?��C�<~�5M��!/a��|��wI���^���z�}�pm�uM�d����<h	q�4�j�:�;�y�!�|����Z�"����
�3�ʅ����T�Y|V��ʮ��<����ūҫ%2��1�
�P'y)�?��c�e�n	�(�����#6eS�H�z��A��S��,s�G�: �[��d�����Jv��"�낃b�>��}��k�V�\�I��»�!�,21ϛRX�wf��'��K$�r��5
��2�l�;א*��C
�8�Ky���ֻ���^HV�N�U�1;��@찖��&P61|���C���eђ�UMlv��C�\l8���^c�]����ё��2��!�h������l8Z�,!A9}�l�p.�w��h�d*�]Y^N�H��f�O��C�k��	��Gag��<����}�qb��q���/�����EU�F{�H#3:6Zb�&�S3w쌣9��2���[V�U3>�n/�
�i�Q
E�VM�W}�������,:x��jY{{Y����;Z��:�zo}���ٺh�F�������9~�4�ZTZ��ঌ����6�=��5G>_�wmQ�8 �ac3�&.=Z�������풐�1�(��Cd�r�R��q7/ )�0�ƁE'�6."J�����s�xǷ����3ħ����K��8ҚI�`�	4��"F{�}Z;3YH�S�,��A��B����0�Q+�Ȱ�(Ȑ
 x��k"�/��w�,��E�8��E\ g!K5$c���4�]m��΄D� ��W�x��`���?*H�U�aш0��-s"�ۖ/��u�>�M�E��f�צq�cI}]d7	��.o�6�J��/���^ّ_j[ i/���7e��=O�M��p��g���ΝR>.�`�g/��R��+ڞ��<�1�Ô/�e)J^C,F2���p���� �$N��d�W��#��cB��ͥ��?�Q������Y���RLЉ�q��~���yh��ش�#$O����Wds�dI�L�8u��n�.�-X0���u�J���3kV�ȅY��uZkC��]��$F�/�}��n��H�|�ۂ�f��id8�팗 �%�h {B��8��@^(�������u�Hƭ���? 밳��݅����{#���-�������JlFS�S�ؾ��)�}�ߵ�Naj�7p�;�.b���3�a��&8�Ba��#G�%��z��޴�8�~��,��>;*���J��*1��ջ$���V�=���v����g���W���Յ�n�"9I����0�U�{���f�tԦ��̲��!�Xm M3RЊJ����}cRo��3mm�ʚ�&�G�
D�����FXi�kޟ@!�Ƣ٥>#�J��g=�u��]a��я5�h>m�_����/�1چ�)�;�d����T��LW/�7�Pc��C<z]��6xI�45�-�	��d�@� A�J"�F�F\B��+�܎�zE�P�sa7S֑��@U�"4��d�l��>�M�D��	���>���T�Ӣ�@x���Q	r�F���w�QnT�~�8Nv@��s�w���'�=F�h�H������U��
�(�T�	H=�f~LY��O���،��i-�O��=�w���s�XՅz�q��y���ߌh�"�:�H��K����8ٌ����1Km{�ǽ�ͤ�*t�@�ߙ.k�ந�	S8��
�J��A����+DJ��f"F��Ėe�aٶ�wڂE���'*�����| ݵ�Zd�K}Jv��HΆ�o���Rņ[t�ð��(W���LJ 2����_���I\���X��2%M	&�?H�κ�1?'��rp�ۇ�TrER���$¢d�U�7�l�]^���;k�����b�L�hLNy�F����{[ V �Y]4g��&6�cpq�m{�0�<E�cdd���A"T�}�6�O ���
�]#Am��޴�x<�O�����3��4�OI_F7��k�U�5�tt>P?ܖz������U����� ���?��0�S���x7|p���\���4�V"�4?p�*�P��H��K�"��?(�Wz�?��ݔ^P8&�Ɂ��c��J�.��l|A,�la�C�v�컃��YG��J��v�Ĺ^�]ktw{�S����OXq�0��y�E���UX�ӧ�ާ��Dz?l���"9�Ǣ�e���,	_k�h�eɎH!�����,�+�����k��oX�+��-z�F��y��Wy.�7M(��Z{Yڒ}���a�w�*���ğ�R���Q@�7wd��H�j�n���5wʉ!�!:��Lt���k"���+5��@��jK��ۋ���~�pvi�`9��o��w��7� ���o9Ӛz
�����O�VB���Rpє��f|x���ܷF��܊���]��*����'�<xaĢ�V����6�]����;��p��W8��[��2��C�䃋���j��+��>�d�?�����Y��	E�"���u�3��f�>`�N!��w�.5�� ��|\\�gl�*�fwE�ߗn�~��Қ8T��àv�����tmGX�`B��rɪ��s�����H���H��zFIЯQ�A@�[6�ד��{p�}En��� A�e6 @�/��xZ�B���R�\od�Ze�c��(!������g��,|�>*q���dh�*�zX��f4�e;�\�3�M(m^oR!p&'cd��Oxe.?-1?/n'��+��yD������O����yR�R��"�e���2pO]hy?�u�*��yTX������@�����1��cZ�|my<�(`MYf�k,���O4@)�g{�I�B#ZE�a��PD$���Zqe��@�>Ӈ���#õ�_.�M߰%Ef7�-����nh���R@p�-�`��y�ܿ�hd�b��,dV(BDu��
���%n�1��E*4�P�T2���x������U
pU���Yxe��M؁�F��C�m�������xO�c 4a�f�q	�f�����!�*��O��_�Ԅ�����|$�9�,0e���)��Lz�J�dYq���e�z�ɪ �����5�4���������Wl�32^��}{����OT�
0����M lT�x@�7⃇�]�� u�[^A+P<,�qa8ֺ38�P��řj����HT��h�$z���P�j��X�L?�0�� %���ள��sc1r�7Mz�=l9�m���k��!�w�_Q�x��r�p���֠���
���sq�.^���&�S��hѳ��x�Zg�]��5�16Xc�β�� f %�0k~6�[�Oj����-��ᬛ&4��n\C��K��n�n/4!X�scT�!/	6�p;X��o��^��[��a,��:����9ao;Lkcp��сs�����qs����uK�p�CL��ƴݹ�W���c�fdB�̳��1�-�VF*T�e�O�v�%�߲����Y�pm��}\�8�x�B�\]N<�pѠ�:=B�5޾'ď�U��3	0��1��`�(�L/#�G�漏����#����l�`��Dގн�3c�h�煏���a7���$[�$�!A�� :U�^!�C^�y� &��p���v��B�I����g�������d񳻗&��]E�k��:�:Ьl9����ߠ�0+��b>��כP�R�g���-sr:ǆצ�p�~<s�;��㣁`k�FW`�1a��Ɋ̈Q��9aV3
�Y�=���Tk�M�6R���J9���˫���n6|��/�h�W~��0�n;`�L�p��=s"Y�������l�~�?[���gN�|E�\�L�N\���C�p���
����c�--��Z�â�ďZ{e�W�CZ4��R�Pi�w��AF<������L�S@kc�[X��.B��`]*aK�~�~^��Kr+yX`�+;n���V.�������?~_"7+n:�v�� *`bd�o�#�+�wlQ����Ee̛����x��^�L�*V�����-��>�
�[/y��
�@�+��4��K��o#��n*��U�w�Bt���륃�ɫ��b����I��A�۪v�[˖1P���(��)mJg���M��y�D@T�ܴ�NBt�E�;U��d'��ZXM��Ǫ.c���7kE�7���cD���c���J��8q5;��X��*�s�Q�kc�@�BN��!k�%p]����]�j ��	�7	�c�0��#�^Xӗ02h���=Ⴂ�wk4���B+�P��*g�@���0�ͨޘ鶻��]�MFbu����A��,��%����şid�Z�� �9��e�
R\e/Սq��]�o��h;1�k� .��O}BQU CZ#��D����x�|�����,�[8E�2r��ѾVֱ��ѫ����q��l -}7�Ϻ�t
�k��7��uݨ�-�����`h���Xi�u�w b}%X[�Z�~=-�BGpZVy$����P�h�?�ú�Mmy�d�Z��Z>M�{��iz5lJ�h~��9��n���ߨ}|�I%=C'��.S�9&�(����i�5)�mJD]���8��L�jT_���CA�X��䈿�7��fp�z���*���ͤ��B��9a ��뢝��B*���~����SI��g屽������V��j!$������z�z0R>�1sC�ю\���y�^1�BTYӡ�JJ���;�F-�98"-'�T� �-~V�-��B�,�Z�s��$�L1Cw`�7@��w�b��\��V6~��D��1���2dC7�8�4fLĕ>F��K���-��&�ƝƼh��٪o�l���6���vpS� �t�AR/�L�-��6@?^�p]8ܟ��1�&st���O����j�J<b~�t}��]X�+��6��m�xU:����S�B:������+�Ƿ�Y���[��B���p�d����@'p�J�t�૛��i�AaRmd�Ϥ�����+R,�I.?B�v��W�-v������B�G�.��l5�}�I.j�E�?ʴ��
�|!rW���q��|���R�m�g�~�u���� �ڨ�I�����â91���J��� j�ś�]k�~�����w����޼[�>�4
��(��:���2[�o�����9t������4�n�dW���D��k��e3���\�� ɬT�h�n�3���%D�n2<�����2_��Ɨ�b�=�P����mV^Tr����V� /}0��	���+H�,y����A����E�ڵ��>�^6(�����~���̺{�Mi��O-�$���L��0�|�����ȜM:�W'��'\��*j�A9��2	�m,�:g�������ʀ����jnK�Z�)�8�_��#+�1I !��ϾaWE������f�!�3+�a����oF��L��������`0~���M&P�ǘ���:���$'w����c��h�F ����-�X�,��X��1��ش�:�h��������_ER���?��R���L�Ǩ�IAJ��p* E�]�h�H��H$-~憐J�/�ζo#���넿8���y�Ћx��g8p �Ρ�A��-iB[ ��}�<��î�K	
im�� �Z�@�,�խ�
W��uG;w({�p���	����9y��'�x�E��h����(a���1M��Tf!X4������("�l�^iC�;f�ߤ��'}x��V$=O��k�+0CJL��aG_���yq7��f4�
��8�
W�g7�Hh�6]f	=[ᒌ�H�-�����%��χI��ո;�Ea� IyG�����ec�>V�����+