XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5D�frؐ���Q��+bp�<�&<�4=�P~�M@��:���`>��q�5����F�Ј���ey����'ws�]�I@�_)�ړn�؂K���J����&a�C�Ef�GQ~��d�4Ӱ�SRAY,���"궇M�6|jaK���^8ƅ�&�q_WSc��:��]w�,�E`��ʟ�w/l�0e�?z�4��[8'��,~���?}���}��X��>�R�shت8�`>Kg|n��\H��3�F>4(d��!�;t������J*5n8�!=z�n�Q�fɞ�^��P�P�q�F�~?e����W���c���|��Ћ=�"�R�H
=s�<,�|�_ˠhI@5q'�b�+j��LJ�{G2�%ѱׁ=�����FJ��[�@����{��i��>���(
�W�#s�Д�]�bL�HE&�<��?/������5@���x�C�E04���*2Vǁ�K��N�0�Nʎ������"�ֻٌ'�*z6]���:�A�_�"p�kz8nm$(�6E�&��,*���7�=ľ�=o�b"��s�!����'�.�&�f����Ĥ �V?�+�4�&gf'��z����@/�t2^39K�Y�K�ү�p��<�X/8�W
={č.��
�Ţ�C�q������r��l�A�PB�N-�u���.���@.�2����_��i�b�)�X�db��y���J�Ǌ���:I��8o���;J��Ěe�1I��:��^|�DlF�n<+p���_}����REH�Am��i�XlxVHYEB    1fc6     b10��V�<���5��f�q�o��u�,�񥜅��絣W��f�Nr[WL~����ק.� ���e|��/ +�����.%��Jo���v%�ߏ�*�czC&����ʷ����?�󜊄��9�<�����LcxZ ��
}�Xv'B�dOE	�(F6�61�1y����zG-7j�"&p��:D�-�����E�tD|�i�7`��	a8>oA䕡�����~���t������̍Z��o� }�D����4p����<<�o=J��m�U-��@iX7��p�@币� �[�/?����S�*���xᶕu�$��D1^ǎw���Hi��GLل�U���b8�v:B�L�aK��S�R籮	���5O[ft������(�R1K�3j���zLi���k�o=��q�̩0�sj�\���GԸ[�6���S��<�tq���`2 vk��h:�ngf횯B}񏦇�C�׫z^���O�E�yK*��=��ӳ�I24�sP��P\�g�6��/*����=��$��ۅ�E/��=������U��*��MQNg�ב��s��~���u2��5�'gT@G�}B��,$��K��q��Վz����'q>+��:Xh�L���3�CCK-.0�?9�Tt��ni�Lp���h��"�A��`1��ϵg$�g������e��D!f���D�q��J�M�QK6�YF/���.B��I�,����/y�F���(v�#�B�����J�S&��x��`���WW �"�hA2!�W�vTx�����̟o�cȈ��`�x}>�H}��F�/v&	���C�1 ��?wg�"����
��Xhcz��Q��1�&��ޙ.�R[d���ȃ8M��}�J���yM����LM�(Ax:�M��	��U	 t�1��F�̣�-M��=d'#)�~w;,�o���Y�j���u�ƍ�υ��C���䚑wYQ'xĒ�J�^��>;.2�פD�H�[�ǏR7%�l�$r5B�S^�?ZG^�Y�
������mh�2O�ON�^;v��#&f�( �Y�ӛ�Ń�+1C�8B�)1k��Y���JG�-��k��	Z2�MV4)c��7G�&���G�i�~?.�^q���v�y?�����H��rÚ$P��Y��3i�`�J|
���k+1������i�S���^4��X�*D�"���b�w�$&����-5�S����֦=Q۰�g�0�MW��p�a�҈�N��t�^��FJYC� b����[ T��b��_��B�9����X5�{Kcq�i����0�K �n��ۓ�Za��7hff�zS]*�I�����ASt�����C�h����X�<�>�4�J�ln��{!��A�wB�Ł��t}Q���8����I�7��rr��2y/=ꁹʲ�=$��*|�]��u��F�z��p��0�rdT?>���d�[�2݄K]gN|-*4��N4e�/^P���	^A��Y
�|!.�ҭ�Sq0Q���L&_���+�|*9Q� �X
�j���g��XqV'�1gː��ܱ�fX)oD��vG�yE������A�����Z�Ӓ���SY���W��O�UnV��3���gI>�6Nu�����ۍ����>�3�X7�9im"2!1	��g�����RW7q���4l|e���h/�f&_TL��h��ڿ���	����!�|گ����z���)����P���_���(�^W�ǘʁ�}��%q?Z��l��~-��qffBr6�$��˜�e9�����?�P>��������IB+�<�*��A�*dnu�_b_u�G���!��b!/�a�5'jp�U
+�ok���V�&3\���RY���`��o��0¡9�Nj�8ν�Y�����v�����4�r�1���oG�>�N��2֖�&x�\�w)���YLT:!����~"��V4В�癰��NH�gG/�>�tF�x����1�_��,ό)|(TB�)W!r~Z�Eےr�q�����a�FL��"i�m㹭|���
{d)�v����qb(��M��U���U�cx��"X����2M��(�ZR�����a�M�Aʺ~+8z6]�<[��lj�{��q�,3y�`> p��Ky��H��%�$׉�&T�0���@F.�xDW�6Wt`��i��`���7.q����}X7�R%W��)"sNn1��*ݾ��$�$�^�c�U|�y(����jAS�_4�	����)^��6�*�Ӵ+mQю��8�����S�=w��7ԖsD�ҧZ쌷]����'�?ny bG����RTWk;��5ew,�87-��8)7�Irq"�aw�O�,1�w1���2�C�Bu��=�m��}�X��w)|#�C���%a�A��G������=34�R@,ʟ������g��zmA�Q{3ׯ��X2/C�!c
�[4*�קw%���3϶��w`��h��5�H�$]�FtԴ��� א �n̒M�n0xTy���/ϯh�j*�!)�}��hxa�x�&Z�x�l.�K�ߐ� f�o����M�2X�B !f�S�'a/WxIut����4���.���iR���Hb�g(��E��yB�H��8V�s��kalWaa>�5L�t�G���niڷ�t��W�v�	+{���kHץEs�V������Px�
��"�R�q2%s��6����U`��Iu�_���Ǜ�8���_lۅ�'.?}�v�[�j��|q&�,Z��.x9��X_Sz����y2�q}�]
���)���)*;@��.va[k���i�q4�!X��