XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$+@nOB���k���Mن�(�b�.��@{Ƌ��)�H�3ȌTʴ�ش,�:�crk��}3����l�V�Hv���ş9@�6��/da���}�����qvE�V�͊x/Bڿ�ɘ�Z���Mp+��X�WL���k-�	+��JZ�;ӡJ�<=&n��g����YٛSr�gN�B;�k9#��ܥ3�߈9�ۖ������u,im�c��H�/��TiН���d$d:������:] \�iJ�:lq-�nA^b�8W�iΛy����W�&) �<���k��k��[w��p¦s�`xt��� -m/S�/���q�S��o9�bP�J��ǔ� ��!�U�v��@��ѭ��щ���o]jـcx��������)m���{Z���6�ĊUA-�bO|�|Y�8�������
���^��0�#�"vg�	�T�bR��P;z&p@n�q5�|;��.O�ޚ������.�Ǎ�Jq��ʦ;N}����1��F����v�(~Z
u��R��S@C���ۙ���:��i�	��e�����^����!��D����������	@J��ڴzoȇG?����l�3��)�����be��&FL��]i�|�-�j�8�B�Ĳw�'����	�L�)��,[rdd��GA�x �*rK���js6#d�=5��� ��V�ޏʨk4���°�n3��#���� �t�˛�] 1��$�b��G���`�G�j��Gg6XlxVHYEB    8afa    1950����q8􁒙g$J� �eC�	���NtR�g-�#��J2�}�Ɛ�4��+s[�9	���ڰ Cɂ�i�K��KXVa��ի$LD7�t��4�Ƙu_��-�:&Ǖ34PU7`�xQ���Tu�FJ6�����(�j��Np>O�Ѯ���Q��ϥ�J�"A���റ���f�RDl׌��fnJB���-����3��$:�jp�!�Qi�A�d��Ё�S�Ǧ��p�(���!�H��U4�Ֆ����]:�����Co4OJ�)%ed�݉�%�@��ؕ�m�<��;EU��LL"�b�L�Q/��ը�ǔ�4�\�`��4��s�^!����
�����?�Z���[�F�]d����`�����D�N��1IV6����HO��eE;���ېψ)�e#�~��,>O����IU'Pr���GWoR�)��*h���)��'�4������6I'6�p��V��,j
���p�u���!�tXI[,oK��߮����#��O[�G���x�d�a�0�ɞ�'>�YMl$��$�ss��-Yɺ����=K'�M�)}�!�{S@���yj@̂q�s/��Qp��I�e�_-�~Rx5�k���!�F?��Z!±�	��-bH���� P��őA�lG��[ч��>���� l��;ϸ��̉���ΔqK�I��ƪ��܅�u?�,HA^�v'��H#?�n7��z�����!IH{"�`xޘ��O��U_�"�I�UrZ
|6vRm�ԫ�SK�: 5y���L$��|ͺ�EB����磤6	p5��
J>t�x��,�R<xqT|�&F������=���c�f����. ��HsK��к7�2�e'zQ`�l��'�xȤF��O�r�}u���߆5p�Uв�^0K9���ܽʅ����?[2�x>��E�_����تFU��R*^��Lp�4u���<*��	D*��j���ی���� �A��)T
�0�z�`���çkr�Aug���_��7���MtkVڛM�P��>�r���RT�y>�Q:3&j��M���`X�&+E�$��2����Ư�""�{�j7|�Z�b-�F������S�]�� 0�)�N�D?�j.n��� BP��Q�Lg��r���O�b8u�.c�l���M�Cꢂez�as�c�?/�|�b�Y���ێ��B�MH:���Κ�ō�?C:�%�N�!��ź�7}�N�(7���_��k#�����2{~���,�sé䛐�X6a��[e�Y�7+�����1�9�H��᠝�l���xH5�B��%�����e.�\�?�ش�ST��zR��B��lhP���ϝڵ�V4��v��/�Ņ1���������P�Ծy>�����c�0���o�k�� ˕kEݞ��s���,���'gh� �����nA��zU������D�wR�!Q�֊3��ؓ/��Н]/[	�$Χs�pѹ�)@��>�7'��jiL���]$i{�D�b���1����lXM��:��gV�B�����D��@	�L�7?����=r��A9]��u�C�����^z�K��;��#��DV�-�)���:���|��c�%�m^��?R�X�m<y���p�-��$��͝�@L/o����a����D�i&|,�hJ;�q�M����a1���m�$Y�V�M�>1l?�>�8JZ�w2�=�0� ���m��J<���<�����:�mk:��.�(Vw���瘰��liF���/��u 3O�w�ͤ'͒_�)9k0��8���O�Ûl���c*Ŀ�Lx��n7��g>`5��G��@��4�Ȍ�T}2�"�~�A>�8
�l�9��"J�G��K3�l2ӕ

���oL|�jN?��ڨa�K3�z��U�%��B���&�PX�?�{e��}H٬nD���]�L�� �0��C+�>��#ڷk҆�=�Z+~6�Yӝ�(v���<���g�ň*���T���+��#� 0O�~��5��a�땄M��w�������ʂkk"���:�4D'.˾Q�R��s9���S��+v@퐺e�9i.��T��n��@�Չ�
��aOD/H�ע�\��Q�B�q6��	J|��$�3U��ґ�bީUܼ�A��I�ǚC����Յ��h����>�$�2f��HW��d�g�G�ߏ��Z�)T/0l+�-��n�;G�W���:�RU�jk��/}އ�J�6������O�̽UhL�����H��s�v>����i���4͑�N�6I9ғ�n���	t�U�_�����������IXE%?�o�ukL��1�i��}=�HP�k�.���P�ɺ���|u/�����<Q����t�@��(���2�p(V�'�'e�,��0�Q{�\�oࡕP�Y ��"Œm��lo�-����[��/�͜VzIx<!5���al�HS�**$:�8�¬����o'%_vU%�
J?0 ����6�U���<Z��d��6�k���g��C���)evdY���G�tB�^�#�`�w}�#I[�ȃ��� ��%,W47�}����H����n�y������=$N�7�s�!؞��Fз2��Ӳ�ӳ��ƾ�f�̡'��".���#�|��ڔrܵ�o���skY���MD�0�_nPr�.��]���@�3Ų7���vi�`�b��*�Divg�f�W}�/�����w�	$����*ƌ�%�i��{v�{0��0��/8����^ܯ^�O�dE��Q�Pm�s�@n���P��Y��^�H�����'E<kQ1#Ly[�;$k�/��I��Z����j�J?]&.���\�H4��8�c+�9��	���������k�V#����T�S��T������S=�J⺤e�ف��# ��E�����8#�/=Y#alI�_v\ ����~��"�aA�z�檯Jb����]m���4�7Л���[,��V� ���8��<�0����ZÅ˲�^͍
�ʎ�N�bV�9a���#r�0D:(�c���ȟJf�m~mz������.w�[�&G���j7sV���9�UAH�
]aG���7����R
[4�����N�bLym*T:���Z6�1+��m�D�!� f���u	�[&�H�zI^B�y�VE�����������y\, �Tvκ ��_2?;6:l-�xK!4z_P*��jq���+�Q�ݾ���]u��ͲW|3��*e ö~j8�<F\\���=�N��$a���f�
���@��M]!br!qu}��6"U����Ώ�GwRV/���?HMa�X���i�Jm��a������7>*y�[dB������n��:S�3�C,9����e�j��4���
(eRYy�����s��BM�#M%��8��CG��~��?�۷��8D^/�a
�~'��^���5�7��hkM\�u��֎f�@gӿ_�3��ti�W��+�O=�Ze���T�zJ����5�9z�*q�Y�H�U�e3��0��)�)�Q��]k��!�U��#z���Fb�O=ȸ�� �p*X����=YaN'��B���סt�w�Q �?ީ1:�Z���̚����{��(�9�<�����u���g�|0�%�n�8&��%�1���
��
k�{xHM�M�_Y�*�����ٙ�L9��UAE-��qQ�'��^�������2H3�mA�6�?�J��C����l-�u˱b��5H�J��lqT�Bi/���i�:�����%L�����+7�U����^%���*e`F�l�� 4�	e1?p����^�'������'�"IϚ�+��M����>�C5���G0GK�(=-Ū�X�����'�6�H؞Q�'fێVi��y6�n��m(|�D��5I,��[���9)���ҵ�����5��jD%Yi*�Z��S��dz��5�,�lA����p��8�<�Q���]��~�=���>L�P&���\,>sU�xe�
��ӆt?��̷q�R*�k�ն&�6+�R���x\��7�{~�g���/���Fɡ�w���ok�m�K��ћ�9�h��ڳ?ړ
�ϻ�+4=���"�����T�!��l�#Кw�:Sv���ݪ�|I�16=��� ��sN���p�1Z���|)�K�JwR�uK}ȓY$�(�L�U7���,��N���jM.�Fz튜CJ����H����nY�ܤ����k/l���U֍�a>캇ɵWx!�7��|�o��5�_=�C{�!'{��5{}�����8�@ 8��XR��c�+h�t���ܼ�s���}W��?�R���uq��6�o�!$a#۩��in��t����r�ᠲ�2)���-<t����=U�R�%m��1�H(�w�\��򆭻!����	�w ��S�h��{D�1�>\2��	� %qu+F�.Ct�*p�[�[�X�u8o�QX
Ow��l��^���@o� np�S��bm�-�%#���'����k�����7?M�㊒�u\�_�%���L %���ӛ��],lf�ceKJj��:X�����֡��Ѐ�-7\nqR���Q��� � �;)��6��6�?��ɹ4��/�R�ұv����;�����?{J�C�y`}�4��ت��LЭ�{˯��a[�Y�O�����A�f�kok0��W,d�^jPsD����m�����ȶ���i���>vpQ�T��u\��}���r��L��}ID���A��V\�H���#�t%������)e:T���^�� I�ҏ�ׯѵ��㼢=��|b/
IJ�����[*2�h:b��1��AB��ڇ�����_�G>{���IJ���%�SL�8t��l�=��,�DI ~$X���O� x��O2��:���<����Q`|���˩��K�y�R����Oi�Fyh��%B��hƊ�)p0�6���,4��o��\����tYB@��0��hYI����y8>|��s�N��u�:hυI8�+�O�V?�t��������g�0J�j��7=�N�2�_ПQ&<�����I��N���J%_��٤]��F�{��Pr�'�#Zς2#F�E3pG7W�������4������3�Rd�@���^�ؤtg�Gͅ]�dWlÖ�G����"��!�\z�ⴜh덓�e��Z��gh=-�����t�k%��l��w,v(Zұ�Mo$�6H�����&;Y�I�_�'2 �a�>�<O=x����yڪ�c:s�^�1F��F�W3h��c wy��sm�\\U�yx ٗ�M��$Ay��\��oD��Uo�GW�����R6b\������](�N��NhiN��f�]%�bBE�k a��U �Ʃ���C�o�Q��Y�Y���.I{���\��4����^Zb��Ky��8Ⱥ��#�(���IP� \��&���=��K眝1�w>��0�E�%��#��T�=ы=0BT�	j�k�?Nf�T��(I�+9.ߵ{:P����?�2��{V�] �~|!� ��>���?:�TF-Jcmv�� J��Ѳ8�H�9�x>%˸����$�����/�b�l�6.�\x���������
 g[��2^���pV
(�j4 �}��0��[
m���e:mo���{ꡌh��:U#Aޓ���L�}#׵�s����0=��9V�/�/���O��g ��|��g {�`��Uz^��s#2$J��� ߫D`J ~o1��s������٪�vjrP4L�|;f1?�N"��촸�ED?� ��6�	DC,�G����GDǍg)�L9�*���h�n���ӈ���������`�+ŏ��_���[�8�/��r�VV�*:� ��VF�Կ'���{=H
�K���ϴ��0�D��:�O���HI�=�Y/`/�T4bx3�G1
�E�}X��wN�Ok�3��3�k��tzxЫ����=:�W11��5�55O���C%�r+U��g���#���u�V|�n4�?����Ǽ:N���o �����AT���'ˮ��#J��`��x/sC{�j�̮�*[��:��cִ�&�р�w�@;+2�fU�F;���7\"8�*��`��yΧ����>&?�����,Vw����8r�e��� &�ϳ�6蚲���I�]۬`e��R3�r@a֐כH<�ų'o �l�7ȓ¡1��ǈ>�g��c�Ǿ��^��(D]d�;<���J/�
�Y"���ia�M�`;�˪�ݺ$�s�ز?�/ )R&��7��$�&����N�N����u�w��'ZMb�-�J��5���V�Z�wI�n��!8L>�u�YL9Sky��������(�A��[wC�����Z�Sc)�r�Q�I(N�0�&�%d���û�:[�=�-���1C@�