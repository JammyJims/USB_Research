XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R��5�0��3ߒ������R�����BE6x1���F����V�vf��]<�#���j"P�4��#j�]j��7w=6�,zKލ��?˷h5���IF�.odg��`�f�����֫*z��	
�I�8�h\U ]���T1v={F�,>��n���(Ed���!w�t��/�~���������-�C"�r2��"��	o�Z��n�'�0S�`lP8�z3��)����X�z�R޶H�����a�WM\�!N+�����Vk�T�Xv4f�gF�3�vn5�G�Hȁ���j�~����ڹ�X��X4'��F����C⯭���tT�N����Y�;�I�e
Z4m�zj#ڭ����������{^�%�w��&;�t��e����i�<&r�J�_��|�ͼ�1]�2k���νD1��>n������~`\�ӥ�/Z/Ό��{{2{]Çn|�{0\t������F�r�m��5�ō>Jy�鐋�g�p���#�},�}Xf�Ya���.�k�v�Ǐ�2H�2��]�v�y�����u{,��Y�`v標-��F�W*� :��d�4�j���C���yD�R=���c�C^X?�/G�P�K\a���3��t5�a�H�}���,�A=?��D��������Z*�w���8s�Z�(T�C����� ��Q׾ьi金.�m�!	��Y��G�������X��4�~�\�0Z��� a��P����W�yd)d%�݇F� ; ۭH�XlxVHYEB    2295     c30��=�+q,
e&0�I|ԣ	�>�Q�K,`��"h�l��j�Q{1%:0$%����_���Y.���PB����h^xF$�&�*f	����2iнY�$U�_���E�zwл��9���z��k�S�T��W-�ל�;d�l%}�v��F
�ed}g'��n�Y"� O�vW��R܀�2�e�ҜJ/G���*�o*Զ���?���^AwU
m'"9��r;���*���)�4Q�m�1�H]�!��N���/tgX�� �/�Z��T��P&Ij�Ll�/�U��^Gp��y�?�O4��w�I�}�gc�Zdқ���1��<���Lئ:d�����E��S�D�f^�hiֆ"���7��r��F-	���ۡ�ݨה5ي�Bc����D�C-��0B�?���3�m��)y�pŲb�i]$"��W�
J�VF���]�N2�^�
1T�����kz�Я�mN���"�}�77��e:_�<����ؐ�u�|�1\��/�Bb�S��>���-�z.nt)+O���dH�`���٣�f�Y.�?-h����%���z�C�1E�r��z�B��>����f�X܌&Sۀ�τ�b��O�礝9�mef�=;jQ���e�'�D���!�^}>�Xt��ٞ˘x��~����Ϛ�P�?��(,w���0?�"e�Ž�+z����
l��g�m(�]��b�D��������p�v�DFI2 ���B���Z��:�*X�%�p�l�Z�Kž�����#�Н�ʋ��C��'S��/�i�SBqf�z����ɒ���ɤ��T=9���'K�ݿ�Q�������z�W�gDli��}��a�����vf�tó��og���Y�\�ߥ���5�c�WA�m�)9֣!�_�$���,�ܖN��/���/�����zK���3
)s�X�OW3�����(-�c*�����0Y�OP��`Z�p7��xv\�1 ��`<sr�|en��?�I��e��WK^�Q%Zh���}�Y�H9�b��di'�F��d`�n�&ߩ}��sJ���H�E�6���˧0]n�ɟ
<]��W�����%�{���̼� S]��sg�]�#���W_g�a��^�x��
Vs���wE�e��2�6r�ի��?]��r�s{��r�źr�%�t�b�D�|�\l�Փ�ϛ����R5)3Y��_���OO!**;�	�(t��d�Y��S?](�87Z��G�B�_�����q�]�FY��!�rqr��� g�($Y-���KW��S�&F�Ʋ ��1���u����<��aH�!�^W�vXc�+���Is��,n�:A�����y6b�x�%�w�w%�ef��򼳀ye�䄤RM�Z�E��Jћ���:�w�#�>�k��I�1���dBF�n:Q����Cw��CHȭsԶ��w�Ԫ?�5�
�S����'��!j���{ӷY9�zU%�Qr���u����m��lk����֕bk�l=��I'�c�&˃��C���H��B��p������DM��В�1�	�%�[�tW��M����<�M��L���@�d�d��᜵�5~#e�H��R���)���_�.pX�]�=��:!�v[,�Q\v�(��^�a[i�c�\�"�J�}������w�?0��V�<��3���Q�Z��s,�\����Z�&X�����E���n�}ݻ<�M'Y^�|U���l�PsܫT�A�;�R����_<V&���r#���������Ba�X1��D��x�e�+�I3G-G��dl)�}��"�   K=�s��jdf4>�Q�r*�?̟��C�I� �A]ƴZ���ݪHU�Dsh�S����i0�J5o�'�&�,�K��/>9B�/i���4 �8��x��0{�F}l�Ѭ�7R�~�W��(��a��ݬ�DH\���L��,ЫB�ph|$_���Ё�� �1fg~h>��@�8�t��)D��<^<jy:tK�-޹ӤG�S#�T��;�b��B�sA�v�L'�s ��_�˫��
Ui1o������:�)
�a<�ua�^�]P�h�rrL`��y��E`Tܾ���@���0�p*ٺ=ʻnY�gV�����_�M�N�	  �9�,+�Dց�V`}�9A�Wٝ����@+h�T~��1=�f����|����PJ�H���5�o�b��1�`��mb8b@G�U4�f���}F}l550A���h��C5ŭ`^鿝����*r9������J�7o-sg����4���fr�����r	<����(�LY2���%.�}�Y"���؍���QK�ɀO�:(���`0�ND�bj�
��x��Z!�,�@��i��K!a�ה>��ĐTȅZ�+���z�t,h����PA���&ͤB��ٮQ��Jf��94U0�%�N�,1��ݠ�Y=�0
Ð�V�sO�{b��>1u����5�!Q�y�S�	֢��Q��8#�`-��ظ�5�����Li$�� k�^�i՜��VH���ܳgxs���&J�/^��rz�s�c�9�}X*Y.š4
{�7R�g�W�� �cQA�4���'4F����<+N�������ate1�Z���L�����gu>gk|�n���s��}���l�č��}��`�Bd�2�a���q���S��mp� �2�'��
��	s�u�M��y�/L.�??�K���~ϓA�e�ɫ�j�zGk�D-���m<���'F5	���5 dx����θ���m�9&v[=��j�Հ�!���X {\=��]Ԇ��u��:�lo��ʼhŖiʘg��-hc�Z�a��RT� �fٔ�
��1����;���U>�V�^��h1�"u>��sn�Pbɘ����|��z(�L6�Ǝ@� p�́�]� �,��(�/i�va��@ c�p��j�>�%%�򟴳A�|*1}4�Ni }Ұ�9���PN��G�^���w�l)�	k�l�uE	�=npHj6�3��P��?�8�xȎ���M
�}E$��@=[h ;g`O_�Q�ԍR=6[@ͤ���C��1!��(���hw��k�@&C�ڍ�
��