XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��XJ|�Nk N�r����D���g���{��.pܢn�'v�-`�+��6�@^���'����x`����R^T�G�Y%�F?/�w)*�K +ֻ�p���a���,nCL���:닔1��kƲP�-��@�u�!Q]����hA-h��5~�`���_��O����XI	R]���&C
=7��5/�G�s`'�K���V���J�ˈ��f>��9dA4�`>m|{�*2��$scdZh�<��Kx���}�y��훞��/O�]����MQ��fTU3؝κ]�p���U�0t�����L��/�H��[n�8�Z��Z�gd�/�]\Z�UA���� k�J�m�Z��֧�N..��t���}��k������}�S/�y�-�"A?-�j��1q���� ^i�S�.���f��Gj���d����D������+�P�Y[Q
�!��j�bK�d�,H���A�ɕ;���^�d�LRLX��J|�4��ɰ�"V\��ٳ�;"هF�[6\�YeK^u���A6����˧X��`=���̻4�9ؓ�o��v��q�R�������9�ks��d�5�5N]1}�n������$�E���eXR;|L3昃�\-Vz)~[f�d�����U~B��{2� -�����&��$NB�`���d�b�"�n����#�kd��}��D���:ɺU}��|�������!N�嶷+r�8aJB�V��PX�j�,~
A�@�~�̴���Gu��h�XlxVHYEB    423c    1350,%*P�p��j���2D+l/2w�[N��r:#w.!��9���~�ӹG5-T}b]�s�����:�T�	p�������R�Ͳ�.^U	����B���^�.Ɗљ:\�}	d���F�Xǰ�E���\e(�J�/F��k~��B�	���7/LK��e�!�F�l$�%{=�����J�4t-��˔l�ƪ_�(�d���2�v}�O��{*�([<��p~���D�[��%��v�*Z,� �OMI�I�2�I_��*��e����F��i��)�z����iq��"5�F/@�,n����D�_B���U''�
z"=�+�E
E�P�f�a�jW^z1$�Vl��箙٧�|�x���+R����ͭ����� �r-J���E�Dn��͘N�K�r��;T�e�Z�7
�9Nr�Wy9�?$��>��3�el9��f��r�W�_
p&Ľ���aj�3��Ob�d��[?�r�5��_,�J�*�Gx��A�ÒG;�@�2���F�K'RP�s:�Xa��u�s��P�(X'c�-e�ڿMe���p8�Dp��C�=�>s�n��ag]/��l:�'��am5r�:f:��+Kbʪ���8���h!b,�7������D0��Rz�m�By���sT��:��k=��b�FlF��g[�GFb�+�Y]w���,'�����w��V�'���dY�+�qپ^^h�BW�����gU��d�d����'s���S�"��e�1W�B6�2m�r��	߶��:,Ԟvp�Dj�h����`��o�X���}`9��!e��/�C�i���:+��W��1IK��F��Z9�[F�:5 �چ]�6B\�V���+��1#���P�s�,�ψ�u��2h�"�l�Y?�tO/F��}�d
��pǹ�%���ٵ�j�g�W&��ĺ"d=�(fV� �2 �}��YT���v���s�q��|�B6q�W�v�Xʏ������t�yǑ�@2���ҋ&K<��󪩛?�ӣe�[�������U��"E0�������� �v-#:��U��s��×7Ut���{�¬����B���k���B��%�	'	j�x�(�M+�%��c�C�����փV����gg� �92h\�<mW��|K�˴�nQ������^���Pۇ� y���
bS(�@9C�/�Y0�8A����p�:��v!
xƂ[pX)���Aܒ���d���KI�z��Y�R%H���u�K2H�+�Y錱��кt'He��˸|<36�JǞ��hdf��*�S��>��VO$Wx�_t�/Ys�_����e�R~��
�m�#�	޴f����8�
���[D���|��"tJ�&*9�t���*� �qk��<g���������7��� ��⼴�9�'��M�@o�ln73�~�Ζ� >s�4�6on݆��#�CN!��$��E�Y��������ؔ}��Z�@"���:$��L�b�q�R��\���,����ʛ��@$��,*A^+���l�YR`0�j����Q��3��k(��lţl;����|��	���U��.�_Mѡ;z��Y�k��� ��1��`����k��X'��\�U���s��^X�Ǒ���+',�{���](��Cj�-�N�/�_=��\�|�f;y�hu���18�qW'_�,�a��/<�n\h_Z������N�Eq[_��dR*�����C�P}�L�}�������'��]P�՜61�d�����/&%��,_�7����گ�s<� 3R�Rf�m�����	R5C��dn�z|��pZ��V7[X�2|�U>���k��zC���v��5��:��/U�t+��o{�1*DB�dF���ǝ��E%W�*!��S�����_l$�����}&T;c����dV˨LF�)��k�7L�ȑ}	���dh*w�췄��o翍��ù��?#��+�+�~��<�-kF{v���'�A��4���͵1w�����@Z�x�G������g�}�]h�^1V��*�m��	�����u}� 㰹����J�14��\ӊ�H7oûq'�f\s��~YF��b�N���ɳHƯ���Қ�U�??fVA�[��U[�/�c�Y�jK���>�ٕ�]*�|�d�/&J�
N�G�1\+U�tzR����[����.�u�P+hR5���5(5�ͬ�3 )��#��>\/W��vZg3���E�8������[p��"��F�ײQvV�3. X������8��K�z�3Cn��'d@�LZ��{�=2���﹡�ց8_�����a���N�G�*�Y�l�x=\z~��a�R�0#-3���d�F�*C҉��\BlK��b+��d'�y�J~B��y��5o�������]n�*�?9����	��qMxg�0��Eg�ĥ/��ך���	�`1D�;�$���l�����'?�(��~/U�T�G�z�d�8���M�[�����+�V��r�%ڜ�[s�Tr�n�+�0���(�y��n��6��<�yPP�AZM)f��8�� �ۏy<8�R��CܛW��Hd6�@yvR_��.6��)C��ڄ�x��},�y��h�+�@N�M�Yh(}�����K=On>F�0P��ɘ�k�֓�/�����K՝�c�6�8��nr�����Q������1�'0��W�X��f�ѡMHV��[�}�!�p��7�+�b�9����q��G�~�7����_�ˁ�du���d���!]Zq<s,��hѨ��ut��ήR�]�[1�TF�Ϟ�`A�X�I��]�W�Eb�b%o����:�Ji����x�ڮg��v�OŴ�x6���1��`U�Ef�(��fA�E@vg��H�6c�%мo�����kQ���IwY��Md^�-lVi6>Rx4�}��=�4��3��,�NN$d����h�r>�l�=�j'[Z�Ne���� �k�(Q���+	#ns��A'�h�F�
c���s4L����YFIl��z4d��zP�yT��6��_Dhx��T�n'����4ݗ�x���>���W4���7ߑ⡃��ֵ�Qd��j�֔3��5�=:r~p�*g0\i𞝡j{�N�+�����i��� U�7�.朢cF�o	=?Sz�	8ނU�vТ.��7#xS#4�-+#`�~*�znһZ�[3'� 
���\�ϘBY��ZX��H&�\vH
L�y��J�^9��ޭNW�J���E5�	[�����\�2����mF~l
^��)ʛt����F�BϬ�s�aR��#�b�13��}>J%sԙܲ4BaL]��^��-O�4>e�e�c-�a˺���
��	�9��$^y�����J$�F���@ g�of�6���,�ɍ���TɌ�I�9}���dʑkўFOwӲJ��[�ޚr�B@{���#���������'G&J+5x�|#���L⁈�� �m(���y�&�:Y0V����M���捼g�\qy���@~���'qGA��zrN�&��~>綘dc�'-Ѭ�_�[/1����HR��Ik�W3�x���y8�E%�Rh��F��(��\؆���0�<P����TԦ�>���+�1�9�4j�q(Һ���7����c��%{�L)�d#�AV��eض̀�զ[ܶ�>Z^bP��R^b�2K���G�ƞ�{Vm�n��K�IY����t*�m�]̟��;�u���٭��]Xm�|�lm��1����"�[Goӽ߁��l�@h����-d��y��6��#��t����he�A�p�X��G�a ΌQ�]�Q�pg[)�D跲i�0��{&�K��"����Q���~�sթ���Pn#Y �K�@y��|�jlM����O��|*��L��V4Ao�Fd�UT��o�;��cc�>ңfR.��T��k����>�D��ƻ���
�j5���b�oUѡ����+����e%�] ����֯as��V�n۸cd����*��N����孅�����Z��
���I��yΟ��������&�'��/t����i�/R�S_�M7�W`��M��[�׫tA8��f,m3k���l��}ɜ{dx(�Hfx9����sZ*���	�8Cd��������"�pӠ���@�ˠa�n%�Q�ɴF�����C�U�)�u%�I?���`5���0��1�|���w��L@}����Q_���	�&���WQ^�d����B󷧝!, �m��Ӣә<�'�N�	?��VE	JD�4F]
ǉ�@�ؖN���Zc�9A<է�B�>;�hΎ��m�-�F5Ut9��(-�JdK��,ŉ:��&y�AD,��rM��3��<��t��e��UB��H/p)`�՜��hp]u���޵����Gq��iRȍ�#be�RH.ݢ`�@�~;N�%�(5���K�_D#IcM��wI��Bc���S�5Xs_3ƒir0�'N��ܐBJ2tZ�򷩰���'k��^�3l��C��V-��B�<VM;�Q���8��ʖ�4�G��U&H0D����`^��������T LN�(c�L K�&g��<Y���+sl�̤�x�^]�rk.�L���;3��Y�Q9�'����"D�G����6
)�N��4?)�Eﭰ:4���R2_w���3._�dwN;!��n(Ə0�-@�S��_m��������+�����W �=�?��B��f����0�v�2�*��}Lg-�A /�L�p+���IX��:_y�W�I�1M5��:"��d 5j��ϭ�l<n�+ËG} b�����V9�%fֿ�Y+N����[�8���T̄�'��_��s��;�j��Xt����.�cKN���R���G�����0�*��R—��X"� �/V��\����8����j�