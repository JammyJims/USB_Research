XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���M��TWX���!��{\Fh3&��I��n`��m0��G9;>[gOÓ���o��]��wI��խ!�+[���t�<�,�n��|��n˜o��_�c��I���m�3����}CG5��xd�=�>��K���k�C�}�T�hDa2{D�*�COd��9����w�g�LP���Yuf�[H$3�KE�E�����/ۆV�)�����
�<���l���(�Lz�	f-���.��em��ٔʡ�/ǧ�~���y�{�-��QI�_
%�=��|X7��=�X�Dw2"����zN���'�h��->��W�$C��]�U�.=��U�-I ]?x?�&�N>i��R~���bc���8����-ƻX�J�_ ��%-�Sކ�?{�Xi�>Vq��teŭY#f���Ƞo��$�3CM~b�*��r� 	�\�}����
g8��}�/��<�yh{x棳�F`>�^7��5�x�P ���{��-������<k�D]:��x���c���Xc��)�L�k�o�_Ƕq��z��;���/g p���R�D� ��[c��ga,!$���a��x3e�@͏�9j4�[��ב �m���IS�1�=�����k�⭎�7���K�B�O�ч�q�Y	̡�,o��{�z�Bo.��B�e��`��D���Z�78/va$ئ�"o*uu�Z# ��cJ�ߢ��6�ZW�o
F��[��S��aJ+ աf[Nt������XlxVHYEB    30ea     df0(���<��(�M큅�AU���u�=��
3r���㿲^<�: Ҳr(�@G	庬�)�Z�pص�8,ij�#�,Un2�c�pMa�5={�a�Nԩ9��׵W��C"�V� ��qbA�@1K_@��0��@��ٞ����v�/��?�{���_�.��9>ҸŨ8�*�-.�Ϋ$Ė=���W D�^�9�|m��S�ω�A3��Z^�xcd�w �Q�U���'���߸��Z��!�쵯�i�|:%T?*Rۈb�"���F}�kݬʂ>�-��]��"��`��Ck���Xsy��� ��vNA;��o/f�j�!�i�>f�e��'V�k��V�K^V��ě��eE�l�6(�9Q ��
&2
n�w�L�����Fn�}�`}ng=x��%G`���Ɓ��֠뤉`QZ����׷NJΟ���XY����ڙ�W�k�H��A��#[��u�<�d�8M^��۳�冾�R[����ĤF�퉅r|�b���<��U5�o����������2z=��4���X�
��A��RyQ�(�t2O-1EK[���/�iK�]
��		�X�W������
��w���}�pz'�WU`��E~�V#w���Y���E��{Z�<�G_��&�6���_�؅��z[a�<��jn]���+QX��Ku�L�K���d�������#�y]V/��ۻn���2ka9i�ӳ�n-����p��M�<�d���I��Y��ꩢNT���ة~ G�"xA[��W�e���o�?I���u�^i摛I�	oڨwvlg�h$�OQ��&����L{1�zhr�u]�-�B3�Lqh�
�VQ�)G������^]`N��,�Z+c������۩��2:{�{J���)~�G��tйH�x����I�`ZE�d��7�����ր��L�HP�+hŌO������/�� �<E	�z��%.r6,N#<�W$��r$�2�|�iJN+,�e��7j��+z�ܤ�zh]u��jY�֪}��8H.�j���G������o<^@���y�?f���lT��ˈ�p"�k��!����.�c�1��P+Jq���მc��������4��SM���<62���ED�$d�<���
pvC��ׯ�8N���jHRMA	�x�+�,�.~�Om���G�Pנ �8w�l�3f�������i1�}5G��R��N��|��G�R4cC�#k|^e��D�K���H����7٬���t�a�z��X=�+qrW���� ꖛ�^�2��N,Xt��Ɣ����պ�/U���\�&��)�0@���眂X�=;�ѓ�s�ϯ��#��DΒ�we)r^qδ�c޺ �����ϣx){a�:Ȋ�om	c�Ӱ��b �P���&fNb�}@�p���c�s��CՆ:Z%*�H�IJ�	�q�Z8�n���������CO-qU����rD�O�V;Ά�A7ݰ+�S�� c  KZ:p�v�Q/m�S��-1 #�m�C�����i��<L3��WR:~�p%�N!S�c�p��$Gl��ŮN6���?�[���
��l�0�=|��b�|oE��E��k��akә4��XW�c6��qƋ�����pր�F����[�Մ��$�-�2v֜V�B�q�?�C.�?\Y<��3w������ŗ	�|s"�t��AOI\\��?�1���3�3��c���W��a�mM���g��4@�;�I��y`M3㥑��(М9(|�ᛜ� ���$���4��xdoh����c���x���v0�ECLO��dօe]�,w�n_1��h����G8�ͻ�~�6M{�/�&k��[�#���l�^�fˈT����у�!�] ��K �"�N�1����7����4g:��(�q����#�l;Z���?��s��p� ���r4%���!P�f���g�l�������9��R^�Z-��O�����oQ���	[�B��tr��|�cWVE���n1���_�8Z�	;�s L/0UhҖ��s|��(��2\�+����>5�b?%�T�u��y��un�.�z[f��$�Y��@b���&��H�Q�PD��:�� ���j��dp����gF�YC�JdE~��&�U	pw��1��b�Aʼ��ͪE���s6p��݅�+���`����l����Gz7+�+E��h,PE�%�w4�΄U���ۜ%�Y0^_��*L�|����;	�5�z�`{��}ŵ����H�de��c<G���[�[g�$���b��/���׋����
��jQ��A�T1�ʿ��@�<�ݍ�S]�!�(]��h;�&�L�Bk)���� ������q�n�bH��v�����rz�_<����N�1��A�kH½3�ԵA�*�3_J��,i��C9z�f/��*�����/��������~�t�S8���<�9s����햢��ʃ�Z�ǈX�-�y�TH�wN���`n����m��d�����E�V�2yt��ZXSXH�)M�"=#���ߗ0�.k�1�w�"^%��qf��H����U���C%܏�4� ��=�Gm7����н�
���V4 z�୻!x�N��d#��L���eWȇ?&Փ�έtLe�Һ��oo�5� pBr�1>�j�4�ͫ�����2z��b]+��w������8��E<6�������l�Q4�A4 ��Y;����#V�P*�-��5��v�C6��]@m�[Q�V�]�4Ft���ca�YםOR�z�{��٤O>u����^�V���NȘ_�(��iڔ�0Z��/��Q���~�2���y��4m�!��\���BK�J��Nݩ�6��6�6�y�n�Gj}�UVY��;A��0����;�>@+�ha�N�R3�
��9q��0��{i���?P�D���M|ݔW����8f|��p����6x</��6��H[d'�h���6B�h��]N���|�)�*�:p����_|�Y�M^����fZ�Nd��o�
$����	>=��`u�
���f?1�	�P׉4�R:8d���L��Y�;�9ov�]�ת�b���w��Ub��)*^A���YP�VN`.b���.���{`=�1�1f��	@m#��Թc6Yb����"+�Xb�����љ���{��@���x-���`�e����C7%JB��i�����M�F��_��;�/�HG����w���JY�]?�$'*˵59���?
�_�xn��%~DoI3�P�M�t?����e3G����/�ܮ,r�^�Yt�׵�E|�����8�T
hde6��j\¥j���m��t��6�}��3O@3�K�`��U�����NWA�T�z}ӵ�����i���AS�/^�I:ue��ܐw��80u%��o��&.o!���,�G����֟��Ag��X�B,�X��/�C��u]�O
��6T�B�������!��
�
c���^�Op>�'����`������+ *|x���o� q��D>��������/(�wA]�5�$��lN��֕��Y�c�+~�u�