XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i�?ZE�b�~-n�BѩF��7��,���/;����R�侃��#�I�$�ng�� �B��Ita�.c]\Γ0�P�u:Jd�9�����&4���p{=��C�8�}>a1��3�Q�OW�uд��*�1�%��n�,]���!u䝬�1�#hI%a�=d}��v���*�b����s���HU'tև�ͼ����Z����c�Ў�Amw��V���ه}�NI��Q�$6��f+��,�A�X�vkY�h�Em�N�݇{��O��oB��a+�EN�AoƋ�x/]�v�O�RC=UY����y��	�%yBy��[/bz9��d<g���U)pC=!�	L�C�/�Z��x}V��iw��m1f�ϽKE�L�^T��y�fV��TJg��M�k��кo�A"w1��)$+�����D�ǧڭ����ϐ@��������mvn��MGWjl�76dBH��<���TX�3��O�Y!
U7CQ=.T�sk�*)
�a�ńb!F�1Y�C/c0�t��r{��HX�j�AĘOLV@�7���n��Byʇ�t|n~k溮�X�m��I	@d�d����m1;��|/�W�B,[O�U���G<�]�5&Sȅm���h����Y��ƕ~�b�9� zoxQ�������ؚ�BW��Uo��>mMe*�����&1ЫoJPa5����o���Nݫ�f����=�����Gk�Q�/�C�BUL���~RZǣޱ�Z��3v��Q>hlV�y�t���]^�\܋�5����c|���JXlxVHYEB    1b3e     4e0���Ռ��bŵ�cYAQ�ZC���Y���@V$Up�N���,n�317٩��4�}��������m ��Qp@���F�%���}3?o�,SR�ʝ�s���[�
�+)�����宯B<OH��ҞV�:�L�s�j��rO��lڤ����9)�s=<%�F�UgL^w	K�?������a�[�1�!���w2�PNV ����S���j�vU1c�:*��`�����|,���V�UtHo�X>���A4��}���o��u��\�`.&��|�"���J�W/Ub7wI)%�W��Xl�v�;�OpIa�f�A�?(w����f�%�6�ѻ������i�/q���T3���˅d�P���b	x�] h�v�~H�׉��q��V!�H���!��å|�T�	E,�;��waJ̭5RD�53U�B�hl&�-����?�[0�y�9��)�m�t�h��R��l���k��NJ/��d�a�ܨ{9������Y����պ����C�
��b�#��Zw��מ ��D����S���Ո�D@to�Ò���X@�M����CI^iyy�B��r%�����ٶ�y���6��a�n|k;��l�����&sQ,o�V�lڹ9G��g�5%��}��!�B` �ӊ��fw�{E��$�)b��NI2m7Ѯ�@
D�.�ќ��?Z��H%3ꐡ���������pj�뺲�ڜ����G�D��.�ei9����aW�r$?���6�˃V��˭h���U(���ܘ���^�Ksj�qu��{�IP{ �F�Kqb}���i���ƮL:�[)�Ȟ֐1D��\���d�<C�pQJ@e���&.�%ɘ ��kpH4�e'6��S��������@3Ւ�)��^�7g�n߶��3|C �-�&Ɉ�S�g�!X�sq`-��.!\���Wz~<�sa����d{SǘO��6�p Q��=3���v��V|�h����r��I)�e��vQo��L'�8���/�n%X���6�'�	���Ubm<)�Uǒ�f�_X'����GI��3�DJM@J|��͢Et����_@�ɩ9��p�#AigJ�ʔɾ	ob�c0I�G��="i@\�wQ��m��M��uj��!��r���A����
wu�FݓrQGgH�!���!�d�[D�;���/4�:�	BL/	r���%貈�_���}��r���\"fea؁��������2���?�"u�_����