XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T���:�T
t�W� 0�9[j��-�Ą��HGGt����#�+�I��=������|[��Z��f/��'!-r5
�^��O���L�~���1T<��Q��W~s�����������Ъ�U�������BcKe����`��Ҋ�13���`���|pu��l�:�۾�Dӧ�����e��9[o���[��N��J&��.E|��Q�b`��/�a&���m�|��yggg�h qF��b@�:�~M*Y�1�M\�`�@hNP����4�����_)xC
���1�9��t���8�.c΄ྒ�Hc�y.�c��wa���bu�m݇ƨ!�E�)W��7�!�/�`e�h���:.1���WΌ ����0�v��i^j�p8o��vd��~i��u��{�m�T�_:�>�)K��q�g��]IU���FL��p�p������`P�_�,�^�Y�(MG��LCU�����	��0�%��JZ7Ⱦ}��a�%S�����䊵-r���Kv��>��]?��8�-�����Z���Y���"P�T<_�t�{a_xE�~�#�OH�?}�҆1����������G��X��*����Y��7n;e,
�\y�m���0پa�zy�lt5����:t���V]v��Z���Hb:a �����H�87G�6�,a�u���<(�\�L�9�v�
��,̌�i�&q�B�.)q��IWa��nB��Z/�{�o�Ku%���I��E'YS��G�"������"����Z��P�suvDs�R�]^XlxVHYEB    4aed    1470�"�|8&��+�R���G�l��_�a�Ob�^~�V��)�v�Q��]^���=��y �
}5φB��5�p��8e���@�;�'m�h�����;vLtB�k7h��U�Ra�� 1�c�,b���&��)�&K�۽�!�p��HY�+5�ô�F��U��#�Xs
x�@��Vtd��.���W&�.Ҫ�{y'�*5��MiU�נ�I0��� V�EC7��Q��J���h9㷸ݠ�|*1P࡯$�rv�6/L҅�Zi/�J:�o�����������E2�C�����J���	w��H�&�Ym}sˊ���5��ⴼ�Z��E���giu�oh��E�h�5'S2���6�������6�C*O�:"*A�-7�~�I
�19H�FEYT�h�.�8bqr&zzOE�3"l�B�qy�Q�F���nLU|;�<�	���)5M	�����G��0�tT2�p[��GO�D��>���Ĉ�롑1����H9��q>/ZC��#�Avs�'{�~�|&��S�O� �"���]|!���'�ʼ"@B�r�o���=|�/ZrΔPf��T5I��� �v�ٱeE�t��5m�"���rzc����$�2h۸)	��1��AT?�QDV�\�䎇ĝ����/}��Mb3�=�ˇhwܻ�%xӜ�P�h��Q�9E�frS���vfg.ɢ�˳�ݭ _�y˴���-P[�Y�3�)��u	8�3t�!-I��Q��uu9V��5����g�n�hO΁薌:U���#��ݠ�vg�e���������IZ���ڴw�fQJ��XC-(^�x]���&���"Z�%ۙ��=�{^a#c�$6Z-	��Rci=�p�l�⎯Ƈv���}��5�����~�eú%��YU��=hkcT�O��0zd�Ƀ�w�_�3����g�V>�����]I���ۮl,�k��B �� �<E9\,#Fz��PX޺Ƚn#��]����tym�_��Dz.S�G�\��ܱ�
C�c�@@��������	-�_$������CсEuＴW�ˣ�v���M��XTS� \��3��o�����T�+����`�-�Н�V�ۓ��̋�T����;^��Z�&L��@d��{���,�X M���l�J�a����A��T�G�"� ᓭϸdX���*�6�����H%��-oa�X�%n�@�ifpn�aV৊�3$�&�����\���Em��(-�;b�u�#�v7�K� J���TV�w�OM͓E��� ��ǋI�C�q!���8(	�ߍ!�KZ�������T�a�2�"{���->��&���O��Nux�R���m^�hE�Oq|J�f���Q&'wּ>��KF���W3��f�gGɾ9S0}ą�AJf�9������ɉ"���V\#�)�)q�B����_�ȟ�>ڙ���"pNg\�8���,��G�a5���l�U�?g�-Þ�[�Wh8�v�β��w'l�WX4�>po� B�U�'�9��[��Y�~���A�����K��p��y1�sb��=��ǯ�����cZ\��EaY4/=�=
�f��I:q
�GD��zT���8��ߡ0ʶ�� ָQ��6^s�g���M�7&����=,x���%��ϲV�\�̱���ri�#���A�������L6G|<�oݢ�"�Xz������a���Qr �M�fKL�O��?�~�N�&5P/Á_|���Gj���ז0�e�� G��j8�i�����сJ���V[t�Ĵg��2j�%�_�-�S��*l|��!�?R�A��OS�,��nD�9��`Ta�m1��]B�+cE4-!�UI��'��+�C��h�� ��_�X��ڏ���ol}��(�z� ��<vT�J�dB��>R���Ѻ��RI�-]g' ��*�Q�GP����0Ѿ�4�����HH��[{��p'��[W�VfK�7j���?�ק��@+;�j��sЏ�-�1~lA��8�g�9�7$�JJ
�}������K�#�{S�vT�_����I�e���đ�����j��d��i���&ZiAkOGif]~(��*[u�0k!���ښRs��Q��Q}�Q�ɉ���I����5���6��E$vs	��W�c�"?�O�O�t��}:-�	���Sc/���<�}L���F�*i#?�n9W�{(K����,�v�QB��."���ar^H|���O�VL/������
xǭ�Cso�>��Z�O�T/�A�{�;   ����1S!^̚�v�Ԭ2 ����FpGJ�p/n���x'R�-�y���]Od�
�~��ZNt��Jev����)l,2|�GP܄R.�����[[H6���w��E�Uɺ��uA@r��r�߭�YF݆��e��BgIl̥ [��H��#��xb�8#��b�����f:�_��4!d��~�ۓ{�ͅ��S�S�%��vt��\[\rm�� �\f��Z+��������
/�y#%n��2<m��b�PV�$���%	�ˈD����X�݆�#c�n���$N�*����"�Y���Y�;:f�}�z�t>���uWsC�Ú�H��YN"�X���$��j7����g
���������̂̇�>݊���ڽ ���k�oH<Q��4H���z�)�B�1��k-��YE��gO�@JN�
�:ksb�˜dm�3r�R����5�t+�e ���3
t�NX���	������,���<��U<A�7�^k'M��hu5���(xAT��q2=Y<yZмe|l����A0�<��v�����H=R�/(O�7�����]%���,S��W�I����P�r�r��� x�@��K��F��ρ%�ݺ���q�I,��x���0I�V2 �jf��3��U/'/Є�q>���u�3���ԡvG��wKٞ�" ��v/*L}��i����b|��O��1cJ[1���5�|��!�*%�X��̞%��5����ykĨ�'N��0��.��%t��k�ݣ���޴Y�RW�^;�;^�l�����)����:�W.�l6ӱa�^@�;26p�7RZ)�o�0(��
�/��V_�M������A0��{��#�p���������5��U6�����~`�]je�eH-r����惝
ɕ����w����ԒD�H�V#;��fcz.�fE}�T���'x"3���-X.	�SY�3�֩�}��W�9|6�m���}C S��b�R;�+��H<}M��&��|κW���x��?�a��cI9��J��h�<ŀ�}���[�q��T�O��5K\�f�?���,C{A��Կ�NP?9�W��6Z,�< *�A�k�(�8Y�Xj��D�I�u�o�\���Ai5�pˈ:n �˙c�"�aOP����Er,�D��8��K�I��aY�#w߿�#��.�^ƕ�|�r�	Oz`���m�%=�^ci�GC�����y�n��5	������/��FN�W��J�"&�:��i�7�t�
�W �(6"��ؙB�Bl�=;�ږ1��3�lm��¨�� ~���}��v���)O�~=Z&��9�;��p����+���ojj*���(g�ߨ�0��j-��\���і�=�f�%_��o�F�of)��u
�9G�G3�ؚ�̭����.Ez���$(sy�m��xL�b�V�(�\Ŀ�������-��F���W���i�E��P,f����࿠F�m�%*�ǿױ܆�ֵy4�X�bV�A�f��@&�|�s��'�y��N?o��@>s��G�)���'���:�:M�L��a���Df���锪ź��}˃r���$hS�5�{��vI�,4�]%��ߨ�r��k��H?�^}��s�^�N������h	���A�2���!_5���.�����ӧR���&#�Y��ؒ���Gqz�fb=�����*>���f�"�'�ܚ�NH���ׂa��);�4��^Ķq ���bs�V�i�H��g9����y�ED<�-��,H��PfHԤ�;��6����ʧ�������A��a\�ݾ������*mG�A���P��ݎ^�%���ʗ&;h���'��#<�|!3i^����s�����;���»��Q��~�F4p�u�{�[��QU;�X��|S��m��@�7s�H�W�'���Qu�}yM�f��֏���"8X�M�L�E����V��7�*ݙ���Y�?[[�r�T-U�\]�{�zUXwb�O�V�;[c�ɐ�]����y�j����f�	9m2
Aϼ 3����u�K����[i�:��{�������OѱC���5Ǒ�c^6�ޯ� 7t�)�U�|��e@��$(Ns���	&�Ei2[8(�|�9���)P�s���x��G��/�`RŃ^k?oI�c���y���K��pذ��4�G峌l/�0�#�@G;e��!����kT;p�.�1i*?�ê�s�!N���+�<7VG��٢ˌp%V=�<�
�ݧ����I��^��$�9�$S�V !�U��2X�54\Y �x�x���g���3��Y���DT��6j*r� 6����Q�7fʃC�K0����r`6�l�B\ȶ��71 �F��ET��Fv�~��v���D���]�-���<ő~$a�	���|hd	���W��Vz<��Y��Qӭ�n������k��?G�l��yj�-�E�l���&Ip���|�Z�fV��0r�Ugt��O(�2�%h*���H�C��dK��o�%r�͟�Y�ᕕi)��\��^���l�"�|~b���(8��'w3�����C�#H��7ǊJ꿡���J��+��f���S����Ԗ.�P�(���8s6[��`��eq0�O)����-��� ��
(2�w��J��R"���Q�i��O.��H{B M)�������FVR�2 �S�~��+�][��r��7��5��7�ac�N@��-�C���=��5�)[���h��U���tx�Y���L�����!��
��?u��\F�Wg���L1���B���ti׶���!��ݓM���&�ڨ��8b�:���Ύ�1�W� H��K)ꡣ.�y!���u���UV�Ǫ|