XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������R�­GJ��0����%�E<�R��gcg0�X���)M�q*��p���iC��~M���\X�ͻi���'L~^vm�0(§��t�T�#Vv�<|L`̬����M��OZ��.�S�[�b�{e�+s�'�B��<�̘�X�5��m�B�]O��k�/���-Q![��";�z������tK@R0��J�.����V������ј_����U�2	�8fa�� �A*b*0:I=�P�� _ҡ7x���ѳ.\����k\Mo��6_�ˢI�(�a�V-q�V�3|�W�tĭT���xC�����"K�r	y�_���m�����FB�����!}Tl��g��w�������yk���k25s*G��P�G���F<;,]�xk�ۯN��cʰ������'q�2�A�Lt�C:f��f���t�-�RN������_�ɟ��H�c9�"��!�/.l�3w˼)�pڄ���,���b�B�e�Ȑ�㽈5g0��ԭЂv�4$pB�g�Akk�B*V?&d�+��G@�����7(�l������Z�����TS��Z�h�P\P�Gb6�`&Kb��{�1���Tl��m���*�&/��0v��O}/�y��'���V�}�0m @��*�]�0���S!z��5��`�r(�ϗ�OE�� G�����͕�q�+��z��^��?sz=7��y�ҡaG��0r�׎���xAw���/d?��%�f�f��$e�K��/ڀ�0��B%�Z𕮊XlxVHYEB    73c4    1220�^�gd@����[7h�;��z���+�VV�7���i�픔hR��^��qH�8���ϫ�q+���	9]f�!B|�"�8�7��ĺŤ��Uʪ圀��#njG�3���@Yj���.-r5���$y��K Y���D�`9��v4�5��镆O)��c�
��@(Q웆�����Y&G#t&�&�4C=��(}����tמ��+�7{c��M����h��s}7�w�x�V�+��x�%�ABͺYqX�Y�R�꣚D�K��C�x�^<P=��=X'U�/�D
��R�����3�c�sv$h�)�ncH�� ���4s��f������j��<�b�'�yp-��.̴X���6'SHV�����'?	ͼ1����ɱ\�~�KD���(�C�o_�\�gLPp�Cw���\S{7+G�(�Ζ��N��K췾D�I�T˧��%�'z��Xa�]Y��6	
{�|6�ŠV�������-�~~�k�+������V$�����̝ �@�g2:D��(�Q����@�S[�6����@}�o�/��y)����t�4b����+��٣��� ��B�k1)	�����v+�y�-�7io��j�uKbG]��	�	tKՏ�{�/���}y�����ǽź�z�
l���9�k��9��LZg�*#��ఐB��� M�n��M�)� y���A��� j���xZ+�5��w��w��E� ;�p��z�wl�(��v�	M��5�.3<]�Q���B�8z?Q�_#�E�h⾝��ׅ�w�e��OfX�0������E���������
b[���ѐ���fI��.a3Æ��?�?����������-���1���C�ҷ�]9&��Nhz�M�y5@g�'�G��0��y�jo�����G����:$�#�qK�w�e����E�����Ϊ/%hq���T�Yqy���]S�p#p��qs�S$���T![�sp`�l�	%_��s����h�v�E���	r �ȏ�\�(|�q��d�Dk�_���@of�4��e�1����@?��<2f� � ��gh��\)Qw��!kܒ�C�6fCDH9�wj����+�i�q�P	]#D]��K}�5�V���\z��r5�2Q�)S���(ϳ��f�{":³ ���vy\4��H��o6p\]7��
��,iϚ�[*ǽ!ZP n~�E:��C96��O��m
��PޭI� ����x��/=_,i�*�Zf��.��G".�P �CK7��ΩR��T,��Px@:/����.�W�j�|��m�:�.���W�'�������L��cmͿӣQ���V���#�L�Vj�wR)�G��ֲ\Q�h�ξ�h�/���,jY�ܓ������A#�����D���G�W���ٗW��
!�wXz?��u�8U�� :GNx�����[������9\RsL��:9�{�y����V�L٪�U"���&p)��[��c����:[��8:�{����c���{��=A�98}!S]!i��Ъd!6���Ԁ�����F`���Q��0ow�k���H]�	F%R��-+�K� ;��ףf�����d��S��MN�~�ziG͞��Q�Y�eщ
����@�Gӑ�=����̺�LH�&���ݨ������E��E��&9���\,�1jPo7ڕ�{刳�Sex�3$y����0��=ҿ�8�:?TS�=d�]+{�e�m,�!;����BB}|1=	R�mӆ���	���ܷƏN(}��1�#^����na�&� �G��A| ʄ`�؊�=�k������W].�ur]���/t�l\[�|+�Saq+0�?$�}��VCo�����n��s�}�=�����1�9���}F�a}��?�}�:��6� �ޮX�n�|�N�.O���CN���d�mCP�RhT�`s ��z.'�i�}o�F>*��JLMr؉��;���fŋH4ㆲaC`.��Y�����l�y�!�6��y�{�*;��ǁ S��g멟���_Ɔm��GC�rA_��������K���(i׷A�L�wɢ^Qy/	�P���[���隴��O�u����QO���R9ք�nw�w���{$����MuT�@f�W>�q���W��rB/k�`5��&eMc��m���9(3��Pcu,�A!���#r�V����I�Z? _�=�Y�����IP�&"��>Ԁ]�Mj�p�KE��.h�GY��¶�s� �Zy4<h�K0�`��f��"�{���S���%B�1|�11��KR!�Až�z����w�l������!^)��K��,�����W=�Y!@$.����3"٣{�j!�QK7�u�:�6ɽ
K��3�BnL���y��;�+��,���78��gM�Zz�����b��U�S��T#�B���,�Z�"�[*��L�o��˄�x��mޏ�Z-Hl���K����f�-H�w���,
�X�]�Z/���������#c�x�(-X���)��c�<���ŀ�A�Uc�:�ZY�t�����0Ր?��[r���X��	Y�8�!�������AP#5D�e�4��G�`��A��NMcSl4U<����n�-t��:.�W�21}RLs��l}��ꋥJ��A��m�Z-���@�J��q���jw87�?CH ^f�=�3���]@�\���j��c<<�؉6�rZy��i�h���������BV����CB�g���-�qL+>[��ODŹXeN��J�f�?ǘ��pU�UL����Pvm����6��PᛎHa���6a�w!��L��[�H-�^qNϚ%�Fz��(,u�Q%�QҲZ�(p��%$��	5.E}k���ejFz¥u�7 -��"�i�qpd�r�Q��Tθ��r���5oF3�n�'�D{�32�K��7i	�Q��x�Z�1P�.���:����_&�/�ڗ�#]S�����P�m|�d�Mk3LN��F����|�t��\h�ў�1"'�0,��9�v�b�.C�q�
�u�5�.xa�ƶ�ɔ�YG3�f�A����0���j���4��gAں�׀�;����w8	���JZ�<bo)�ڃs�#y^q�o~W��}bh�T��-�}.�l_g��R0�-h��}f���}{Yؽ�U�jM'˶�y|f3��	C�)�um�*Pig:Ͼ}2Ғn������� ��y<f���B�,��|ԁ�K6/vR�0�"x9"�}6�	FD�d���s����4���I��M
ʘ�������\Wo:Sy����9$ ;�Hnt�0��$�r/L6�揂^Hy�}�~ȑr�B��1�$��2����f��	��
���ގ�>��R7 �te�����6��ˋ�xYk��0Mkd.�R�r��BNC�D����>X0��rsk*l���Xwd��$_����3(�[l�
��a�,Ж��ƔH*<!ZF�xN�A>PJ#ij��aBh��G�U࣯�YC|���d:U�(�/Ψ))Sţ���G���;�������]���h+o^D?^��G	�����ׯ"�Vzd�W�,�Z#�y�|��^�8��}���� -{`p0oj�U�WQ�Ld�4���C�����W/�%��2��ԭ��e�yp[���U��T.zy�V�{��]8�b��[��k8e����:�]�k�E�Hm0��7�y��6�y@�2b�v+�=q���K�0c��!��v$`�4_��~qSW��N��{}=677�l�3I�@!)v/�t �A�y�cû�_�O���� uFr`�9�=<{{g�Ѓ��^���4 |WJ�C(�O{�����3�dm�苃�I�Z^�1e�Z�RR1�(�&�{��2�Уv�+�R�m��=�Qy��
�g^��=�ZvS�X�ӷ�cg?+���>���D��k��M�Bw�gt����������֪�P�'LDI�//=�)Ptn�Ԣ=~��0��S@��>��|���@L��?4��KN����x*�������%'�|�&��:�w/�4̌8��^��i����(�vO�Dò~��W~Y�H���ک�K�tzq��P4Nz̶g-�d�1��m suI_Z��p��8�'](��$�����d-_P1��~
SJ7�-ğ����s�-Z�?)���%q�OԨt�,A���	�f��h�]�sQ/�@_��+d�>!e@Yl�����_����I���>�*-�����Ƶʰ1�3H��Ĵoj^RO�v׹���f�˺瞋�5):(���[K�˽4��4���4$�Pi"�mȘ�̻�O 	��;�s�/�v�xo ����S���̩&8���7|�W��D蹢>pb��;?��8��*4��T9D�B_1�l��wC:'nS�I�<Qm��<o�n�����(��A��3^{ԶM���h	S��b�|AZ�1������q|
�F��ۅ�ip��|	WC �|[@�b"�)���P:+�d��lJ���A�jA�~����g�}�+� �bF���9����;:�^�{�K{>,v�r��%V�pc�Q�ެ2s���S��2��ٖ�u���.~v��8�c�����n"���mT�U���Dͥ�2�=