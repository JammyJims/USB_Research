XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���x���ՌI���@������3	s����ɽ;���o�f�H�x��伯S�@R(�	�Ü�|8��a���y�7�"��B��Ԇ��"�#����=k������N�wh�GR���Η�`�sU���\���s, �{iU7���,���l�p1��$C�iN�2E�j6,����ޠ·�%�!r����! ���*���>��5)0#Oj-��v�������i�!�A޳z�_io������+��LÝ��O�d��gWY�m�n�p
I��($x)�j� ��t�0��欜`D5$��E����h�1�T�ńy RdC7*O�ي��`2R�*J�;�������3,��)[�!&�l{(��t@�=�}Ĺ&��:\�9_��5�˽J4�{�V��x@��&���ť|�;|��RO,6d<B(~E�[��I�C��a+Y�o�dk7ݍ2�<���bl>~��q�����b��e�b"�1!P�-�4�b[$I�y��
"�T�/�A���hZ >�_`���LB���]�^�%�������[J2}s-;U����(�4j�>ì"��7�EGA��4׳���<O؄��^�B�1��2x�{��p���^{%rQOu�6����� j�CR<��#�"�����m$9Cp�'��Y;�v]e�׏�"Ǭ]�T�7�ʡ:�?��(��y�/u�&�u��Z?w���8�sᰙ�ť����
]�ڳ�15fP�=2�T�&7E��Ƶ�!m��{�����ZXlxVHYEB    22f5     a60e���6CT�-�|��lԼ���M,�7�"����8�*tv�[/��!��9��9F���Q�S��z��\l5ѳJxY�����q���9oĔ>P�LP�G:�B�|= ��t��Eq7��s�"'�W���� :^� 4{(�X�Xgʌีd�9���Xs�C�O�X�A9Lo����w�mQ?��Q�d��F+$�O7����}��e"�X��@����ݨN*��K�\i����k$�aY��Ú)SdܢC6h��/pĶ|Tغ��)�(j[���ofS:�S��'�9�p����� 	�T����{�~r[���]���=90S��i�4�U9R�q�����CDO�Väcw���d�6�d��gv*�� "�ZIZ�Ƴ���	����6K�K<KH��ɀa'�w	�	k��1̮єUv��λ��!�<� p��b�Q�Ε �ي�5���Sg6`���y���KU�V�2�=�0��þ�z\Tn�0�}5�3���83D�D�������g�;�/�ΐ�jW,YV&�j�󢗭gyj��#�t�E�ꎳ��4\�Nx]��e�X�ԭ)�W]%u�
|`Pv����Q���
��I��9��ڣ�~�VΖ����H�3����HΟu�EE��JB���:�hy��=!IXi�8V"O[����+m�ό��D����h�s�t��-��<�D��Z�
;s��Gos����V	�����Z�=u��ne�2o� ���!qށ�����t?X�E���"!U��x�-�O�����,'��rP.1��B�_uX�Q�j�a� H|>ú���?��W���Y��(���D[~��(s�GДT�,}|�&R'�&�o��uwz��7��t JUe�D��f�xe�'��mu&��� ���m��Η�����v��.�S��E���Y�T>A��Ȑf�H1�,��}���Ő���qG�<pK�n��l��EA�����쑢g��׵U�.Fa�&������*��n�_*���uMH@��K�.n�s���� �(2
�7��Z=>�h+��_烸~p��N=�X���©O��~5��!Y)�*#��W���O|e^�b�کމ�O���#V���,���c�w����"U���O��*��Au�2�N1���d��ٻ�E9�$\=8&5����0��WA54��dE�_zAz�pU�H�Wgi]*��K�4O�Cж������O� 2G6���	���WZVNz.�(`�[�v�p�3�T�6��J����e��.o���uq
2�]�SY�{.W�+���1��'Az� 4ݩ�%Ts�r��l��~ }�w��~��=w�'���\�l��)��+�����f��Uw��~�05���HF0�/�Z?��n4W��U=z|5��e��֏�kZ���m�`#������J�6#2,<U<qO������ށ������ܚ.f�$=(�yh�rf��:/+��}�Y��~��o={��M[�h7�jm
��ym��5ٴ 4!��V��	�Z���hc��h���	�y�R��᛬0T�Jx�}���)��#���|�F3y���l`#�+�	�LC����[�/D��\ʬ �
��W}C/{C�!��n+ �X�'�"cb��p�S�R8×C�Ư��.���Ճ5˝W��);�K��D2�SC�8XaKD�[����8K��:[m�ñ���fXU׵#��{N&�9��NӍ@�0�+��Aܤ֠���4��ۼދL0��S*b������:�c�=���@dl^����F�����;����!����r�O�F��EV�,+�V%��Sh�>�yI�_��K��2C��!��rvqo�W�6*�ߤSl�H���_�
8mϥω����g�3�l��D���S��V�Ƭ^a��N�5
�:w������`<�e�E�@��J�$�?�O;�������9���כО��|��O��h��Me����P�`�!k���E��H	^�O��($a#�p.H��MΑ������Zߖ���$!XFߟ[.�#�e�"f��N�D@����=�	���쉂� C�v��v5+,^~$�Mz,�V���מ�D���%�O(zݓ��~1�ɯF�5Uh+�
�x���+g�~�E�8m����8��aw�S5����#N�ǹg�������Ȓ���s�mt%WӼ{"ye1!���S����V����b�'ãv(��(R:^,u]�|��;@<��9VU����m%�D(�i���C�p�����d�[e|��b[��z���8n�OIw�ޅaJ�V�����1p���g�>�4aވҼ
4!�K������(�ay�p}�㢁1'��P�����]�M���RoJp�l;E6�qg�ϡ���-�L0�,����g�H�?.9��g�D�����d���JOObr�A9�=Qr��+c�p��\n�>T�j,O
{B�Z�f�r?4���T��>��L�.���P�/*	X�b{9܀.�����F�>��J���������$-�t�k�$��fvM"9^�8�<Ob����N�5��Ǔp0	�I3��<,ƛf��gϦa�B��܋�P�ߠ%G�>
��l��cNRq��~�5�[`�