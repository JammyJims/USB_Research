XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X��C�j瓬j���"�p�۟eR�A\ͫ%��!@�@�ثfv�:d�|�`
� ��s��扺t� ��Q��&��Z$Y5
K#����Q��]4��
T�6 �G	i�]i��d��~M����H��.Нt�J{R=���U�K��C����5�I��A�Bs��N�°�-�� �j��#��
�!}E (A_�Mļ�Y� DRˬ<����N��@����H�>���'��9���Q[8�{�D��7ALJ�2TJ��T��V:����]��.�r����E[c,�ݒۦ=گ���Oh .�%-�E�_�63�b?����is��i��G
a���&�X9�Kb~�{!��7��ل�05�- 2��ˊ|��	g����Y�y�C�n7E}to|����%HuJ)6���,#���<�?��R��Z���2\+�1��?��7o��C���.}Q�x-����B�c=����hV4��9���N\�٢%Z�|2r�x�ȧ"2+u�Gv۹��¾�ʫ��at͵�����
��e;�{���	z
+�2(�SX��k5މ�k)�CKJ?�[/��B�/�׀�l�[Q�ZH��7�wa�Z~�����b?��-�~hH���+_\��ex���p�r�\;�����.���8�3� N��6N!�า�����
�jٹ��)�W֟��qndϨWWf:�X�k�9n�������Hv�t��ëd�8U�XD��[QQ`�D7c��6�*���	��XlxVHYEB    fa00    2370��^�0$X�M1���F�c�,�?�Q^Y`�e*�� ~��Q��ս(P	r~�L��b�O`�Pm�A��K�#\���ԃ4>��'�Y��ދU��"�_�,ϳ��~�	tg�(���C�	��C�;j����������.6
i������8�GwD���3T��xe~)�����uH}2����\�#�U��Q*�4%�A㍹N�m|��]���d����9�l3si���aѦaN-K"솺]W����YhZ�^<�TLa i��iw��"�s4U�6T�S�R���2ɾ�1�Vx���e1�<�1��W����\."��X�ŀ�m�$��3S�pk�h�-�S�]?���a[�N��>;I�_]|I��Q�4����"�?���.ʙžO�$�3���M��V��������(l��"���R�6'F����A4��	P��#�R�	�/$��cn�*}f��3��$����ᵚq4�Wn@)��g"e�>�5�x�3H�4�x|�t�q������
3���>��ϖȬAX7�QpvE2�'�Op���8w�,�y��A���Pʰ�INj��y���s�d�}�G�N����"�# ג�|��F�Li��N[B�BD6����51����^Z^�6f�K&�� UԷ�굃|�	x�=�绋|��{\���c5w�Y��ZtCj�$X}y".�n��P>q�B,�nj���$�p���R�H����;"���}pg�q7,�?��$	�&��
���CI��~���[�4Ц#}|��}tx�i�^j�F�]�2dF��r��SZ%���Eh*���6)dx�5�4������/��>���S��)Z�i�z�]������!��|�d/�퀃9��w��5��)���bLG����7~�T�+cUG�3�҂����&�]怀�&���ɵ��?ʭ��͟�׷(�<�UH�>_���	]ڼ���jye��g��¡�C����4�m��8Xժ�U��(��J�<а@�������$�6b�"�s�|H9�i�w�N��n.Ԝȅ!;�k�
��y�l�p�������L?����3n�>�[V�f���]�u�8G��n�ͲC�M�{Цw�hq���t%W��9�o;
5�З�c�Z�Ë[$¯����E�� �V-*�1���À8�Ue��t��Շ��n�{'=�+v�d��J�����x��}R�KW:֌��A��D/��[P�fݹ�r�������E�����oi�614n�{l8�u��M�BS��7Y�3iYe��zU���S�7�����)oρ�9z춌C��2s2��-���ڧ�P�^�1�PH�OK	�>XX�m00� 	*3�)���ce ��+&��,����A8�2<pJ��V�F_��i�&�Whk+�E~���|�ɟ��r��5
(�5���,"�$7�����.�в?#���Ⱥ-0t@3�p$xp_���*���0��Z�'��"͇�z����������҉5�o)&��H+z�u�П�� Ն�~15ӓSb��=���:�2�Z�� �>�v!�ҳ���jzT���Pu ݶ�����[����yipH[i��MNjgco��`h�O��..XDm6�m�F���jc����g�>f�;�
��@١ᤚ�I�x'��z�ǘ%�}�5o��bZ���1g�eO�IFT� |T�A �F��_��G�{+��@�t�՞@5�{[������.1�!��P���,�Q��lˮ��y��m��>d��ж�0���s�t�Rg�X[��~5,!���럊�"es���6\1�����D^��w��ͧ�S(�AfL�*�@��"��uTU�9q���X�܂J�F!��ƈ��f�-�S��۞Y��'�����IB����2a]oi�4k��&�Jt�ٻ��|� �Y_��i[��E��z'd�\w��cV5�S�C�03�^,L+l�}��n�/�39<6���U��c��Ƞ��G�2$x��ú�y�`M�U���CJ���1ζ�1_��l��7�F.h���`���\_���!&MO;��A�x��ϯ���'9PD�]�6�;;5���;��_T�݃/dr����U^��ʓ�s�>��#gK�&�ϑ��h��}�ԻA���6� ��F^�u��֝�fD�4j��C\y#�A�U1E$eJ���x3���,V�\��>���l�h'a3g����hV0�K��8ׅ��-�����t%{M�q�O|V�0���=x���Ủ��oe�f���ɘ�)p���9VT���pG>�Z�^��4��"T��)Z��sg�՗���-�G�s���}�n"20:d��aق�c�}�%�f� �n'K�����
��	;%� @q��R[7�Nn�h�%��G��8�y9��{'4S#�X2��"�\�����$�)��E}�'M�8������ٓ�w]�]�}�U�}���)R�d���h�}Ѻ�${d�N��]S�`{����r��1n�斒;o4��ꉂ#�T�yN��.Z�1��dTu��;�_���c�m�+����j.�z��ʲ���g��w��wQ���C���ЊR|=��=�`���.�S{gsQ^��]y����I>Hb9νPu�u2[�w�^������Q�$��Rq"�<ds�����dy��d�f��|E���h x��#o�����*׏dg��Hk#�Ag]w�C~0.{���;� ��ȊfE�d��\��q
��Ĵւ��И���k; %[i���z֥��w_�}��� �9G'YR�
k��h��η���Y7$k]WAr)IG����]�v��6	������j�rJY��[���BfN�����k��#�bʳ��� FG�Ќ׼�4���i���in��ws�c�8TzJ� �+ɳ���翶�]dXLy���@���3�I�?Y�����
�j�����B�Xb�!]�杍 7�����vD1WD�=���t�cf��G�j���-��l���-����4����y&1�4/����cڵ!�No�qz�!ث�"�t#�eҤ�U�A�rv
�\���O��:��Ip����v��aK3�scABo~i��7��΃i�6�Ium��4}��y�uM0},D�4_��@��OsԬ�swC�7�,��#�S����S�N��ɼ�vގb��j���)�]g�%s�j#ca�*�rϘ��T��[U�\�0�z�>\���3:$L4}�L���%�_�@� �+�n�D���o�Ax(=Y�X�%X�v&梅�r(�����>)!�y3�5���ڀ�|М���MI�?16��%���N-�� ���?3�G�c�`����,;�OPU���
;Ŀ���ZlOva�L��ǻW�����*��q`��8��{x��F&�$�G���&�q�]&2ޘ- �Ҏ�XC��Oz���8
b�N�Dw����Fܦ�Z]�ؠ��D�C<q����}��P 4�*�e#�᫚����kq�Q������@�&A�3� .�|�a�N�R�Ex����v�-�c.W(!"_2�u��~�?P�-!�Yй��=1��c�HY:��0h�E�ԠA�*�ݰ�6؂�$�;���ڻLu���@�<��Z!�_p���jT:?�p��)�����+��K)��!���+�I��֛[v���&�V`�d�.H��9�Cyr��#r���Х97ԒI/�;�kEC��@�z��X�%0h�@�iꔐi?m�_x�m"#��fZ�(�"��\)��uϰ����m�wg�jC��w�����%r�lf���};��l�M@������BE���ٽ�k��@�����P~�z�G�D���~:$I�g�wS?��{n���0����n*�!r�~���9o�nG3b�������}7S-"�<��|�8�F� �	W[+��-�>c�<�X�ަ`���g<4�i����
����*����Fvh�f��T��:fi��Ӈ��8�'P���"5�-x�D|����?Y.�>V#6���"���%�d����o��U�v�*u	4�Z� �&;įP�ؔ���"�2�<�W �2�����o�!hͅ���4�>s'&u�^aՊQ�d���{�,�SP]�E�]��}1���&�F���o��5�'x��Iڜ�%�ŏ�0�qq�ՙ��\Q3p���g�͚Ժ|�F�e[L F�¦�K��8����:X]�UлF���1�n"��գ����D�n�]�C�'��.�\#VP���}���/7\�:DDU�õ��{Ɉ�:d�p	�y,�����oT��A��N��{�e�r(6�|@���.�#ƶؗ�(�%K��h�7�L��-K����N����1_0vΏi�xwT`�c��S�@럇J�c	u�$���l���7�M�kP��;�-u\BDc^�3)��	�|/�oF�����m�@�j�e��/���W�t4�?�x���>u����Ǹ��u94�g�QH��ܵ+��E�nt�X:��u�)�@����C�g�6.�!�`!R�Vg6���J|�!���]�"Z��=�{�'s~�/��F���2� �LBb���';V��+kA�0�v�(�,�]R���̣r1��
w�5L�&|=�M����6��(�w;����g�-!���]ދb\C!F����38<>���G����tZ�����xb��H�Ҫ����G�V7��b C�:�<�X��ǾC�|Ҫ\׏����Fې_!tw�>2j�Wr��C�� �7��{�����c�ٲlv�B*w3�,�b�*~^Œ�z(�'����oJ�����CTD���Up&�uޥV剆G1�3������lJ�'�i6��'(��n�2�5"��:�4=�/N�&YF�q!�X:�z�E��a��z1���e98���}Q��a�ڂ���
��M+>r���\��H���28 v���V��� �e��`B�k]���U'�Wq���Uޫ.e|6^�t����zH~���	�R��Y)��LXY�ɪy�h�ܔe�`֯��A�ab�Ex��l��-�5�L�(j�5:���1}CCX��`�~�M_co��K�mI[�u���zGԔ��\.Ǐ�A7'��df
S�����]��wt�G�~�N܁�?`��x����ed1m���}��h��
�֭D49����==����|Į�t,/�/OYp{
/�$AN�� �����M���*

��]6��`��ʟCB05	(ogu��G���T�z����@��s�sq'�ľyb���;�E�Tڧ�hc^I�n�c��+��>�ד𤴌_Xg�I���q�U�w���K��|�e"�y2A��3OJd4�<��@4Nv�3���5�^�_��i[B�F��a�$�m�<woi�/\���7� ���vb
qq
�څ�],j}��8�?[��h�p���߹w�=#3/��� vt#�Y��n�V#�@�0�1�;���N
��nv)B<#_'�ӕ4�2O�8�1��xoܼkY�!�?�V�/�!Rї
��tk��66r����Ȁ������)�1&��:��p)8t{�4�� ʀ9/�����%�%�3Q(;B5��X������(˟o�;c+ܹ䠶�_����%B���9�T�'�S&�X��;��Æ1�] ��Ĵ�ݞ����5�~�ZJ��ae�;mQ���g�(��ȴ�u��$�
C�ƺw���@Y]�!�������ϔFzV�K~"�T��,X M��r���h����ߝ�d�
��Wb��r���7VX��Në�"��?SY�ps��Z��7���C�<%F	�E-b#�9��{���%b�uh\��������t`lZ��H�h�g����{�Bw3�_� �:/�:\�C�����0>Cf�͎��Eߦ�}�7 /u>��Bs, �q�U��V����ohk<��eo@%�;:�x���Vxzt\ji�#B������E-���6�N$��g!�:��ٿ��fi���Y��H��W=��RTD��'�H�y�*1yH�W��a�5�E�UP�y\T�������n��mʰ����s�Cz'�.Ґ<�>Yf��1��?�+�U!��(��C��.y�!�tr�ӕBY�_|JY�L7_�g�pFO��6:@C��h\�L���������U�� T�o~g�g��\����H:+�g���Rq0��\c�Y����TI<}���=�s�7��wI��V��`�HU��o_�s����g==��#�g�:,ܫ�$>�������T��ψmFf�g}�۾&]Q�]��EG@�]j�C�mr�"��'����] DCPj�ws�-��:(�ig`6|"�S�z8�1�p�w������*�y��p�d_��`kD�JKH;0Ďni:vg�R��I�[��ʸ���#�ؠ�qC�)"��̫5���P!��:gdP��l���I���
���ͭ51�,j[���º.���,�1�n�D��~���(�Q=U������H�nk꿧ʊ�<�8�cx�ë��\u����')C��Z�v��z�m�1�����m)Dw�t�R8�p	�Mm5i7�a��>�>7��	��x7���S�$�R���҉�4އq���Z"���meq=�.Q�U2.��oB,�K)�*8"h�d���c�������}��U��)�6�)�-�p�Y>�Cߦ%i|'�����wh#ݯ��u-�n�aQ������n4$lR���dW�;�X��7M��W��mrհ^���܎��Z�5u4�=I�b7�<���Ň��Uh�cuc��$���mbL�413�F"k1qO�lJ\F�r����+�2��c`�"���/�\�jcr�%Y$spC�l�$F{NWm��]6	�t�V�"��s��)��P��3`A���5����0b�eGN���3:�_Z��[u��[8h�0�uy����P'o�c����2���\x�*�	9 ���2�B����2idL�`?��j�6�	�8O�}8 ��0�mn/��HsQ����Nze����A�V�qf��p�2y��j����Oj/�օ��Ҵ �>X�7!��Iub���gI�%jC�M&/��E���f��|���w�	�π@����.'
�OX����1PFP��>���`I�6�F���4�x�6�?:H�k2\e`��8w�'���s�?�_(n���+rQT1��
����Ÿ��������ܮX5��б�j�!L�b���Y&&�������$7l � 
5+�7�C�s��/R�C�����ձ:�u�4���kHQ�A�4?����GD-Tr:� bC!�+�kml[�eO�N=3�$�R1��tnb�x�}�.-�[;g`��7�|���-�F��t�V8�R�Y�{���������e��N۟bd��oҍ~.�
G6O�e����3�}b�X�|�t�X"��P����v�3��t�n�+���8��Е0y�a[�x���Ƽ��XMI�ϮK�>�K�r+���14�+�{_Rt���P&ۄ �c�iV���".��;sRaI�>W����wHy�H�s~쏔�[fT%$��z^��C��������W�b�i�R�)L��;�0J ������A3yN��V5l� B8�9y�&�W<&�FY�,�� �n����B�a���C�\R9�}�
�1 �;r�曐4_�&N�*ƅ�o�U�g4�/6Jv�ج��ae��C�;�H����ws�"�O��rtK@��,֨e��]�z���Fd�@���&��r�Λ f9�F!�1 e�<PG�3�A�s��!�D']� �&��,缑��̏��Y�)-��e-'��P�����R��U`
h~�ގ醁�0Q����-����T�I7�[�Ej�L�����@��&��C/��{Yj8��o�u���AI$-��!hۛ�?_X�ˌ]�̪�1�|���|���������x��{\7lكݨ�*}j�|��ル�I�X�z�
��t���z"���� �(���@L��lj�hZ^TɡΧc�����1U����!�V�*��o$ş�^�C�[����L2���j�tG�� �{6q����G7��'P�W��8c72$�_���ԏu
H��3�#q�ӫ�%�f��m!�� �3���'�uw�'$J�׌�V�����A5x�1Q���j�x/�kf����,�a��t㻚*A
��Y�����la����mS)Q�t�\��8���8'a'l�K���a;g>�6�ab?�n0���XV��OߊB��8W�4f�g.Q?��D�͌�ujhZ����s)�̼IV���y�k�4�>-
����o�~"�F!SKE��̍HW`Q�E)��g�}@�����"����`=��$YQ���ՉN��ݜ��^CQE:%��r�����Ύ,:^ŕيu
=|��]}�P���W}���b쯯�9)q!a	!k�Gg�,��A���\�"s��r<єeJ�/?p���P�£:�@?�"�p�@f�Ɂ��>�;h�}j�)�mW;2{�/�y�J���P�ظ8	����}:l�k��C>����9�C\����Z�Ւ��YR<6D]���8�Lwj�4���l|`�f�X,`��0��d����~ѫ�
�$]cڢ{��Rc��&��;�2�����j v���V��~�MB_���U?մ���}�I�5n���)D�M���O߫���6\h���1=S��,RՋ�Z�hMCh|Ư<��,�8�l���M��HY��Y� �e:�#�~%�}��o�s5u�3�jB�/8V
��e��I��+�O��ss
��IR�,͟���T/wT����m�d�b!��ƪ�e 63�G�	���d1n�r�a��n�z��2�Af�4~��o�ظ��4?��y�߷�lٜX�F�iH_1�R�7_����T,$Q�Lq;������S��e�)(ь	])_���@�⺨b*D�6�����x�Q~b}��푤�݋���Y{�y1#;���&Lфn����v��XlxVHYEB    fa00    1160ygsl�W�<�l��F!['�V���EKH�H�ޱ������Y�+1��Ҧj��Փw���H: [4�Q��B�#/��P�nb�s���(�����TJq��SZd�#25�/�JL��M�����67������2�3�`�����b�,�����0#��ۛ����_���c�c�| h����E�e�,�|v�J��PՎ	�\ �G�9� o��A�z�E)t����PnUV��l�3*h)UD�3��Cب���f�i�-�o�e/��������3X���nQ����m�&�q%*����/yS�H�k��6�֣��2���2�L��>�58��6$� Zr�"��/v�J����	7�{�ґ5&��\j΃,F�:�Ŝ�ڷ��G8�P^�3˪4_`�P@Zg[�:d��������M͘��׸='�B_��P����L�57f9�"1º�V�ٿdt�A_�KN;�6f�TAbI�T�>[�<�P��y��}n lݜ㈮�Y�E�eh�V�n>��nT������s9��D���f�'CCre:�5*�����%��q�WB4h�w;���G�[u�e���ug�q[|�dɱ��ݞ��,f>�3���2ĐE�@N�/�'SRS�/�^�Z$ɐ��	�� ��!P�ПK~Q]c� [��NR�[K"J�W�	�i`�W�f��{R�|(X!k৓�[�Cǁ'a2����x���!�uI3�N�i�����]�f�%^z��(�i�k����������Rڕo��REs��ȯz��y����(�Ym�n�kC��ȿ����b}N��7�a���h�Y<{��d���f�e���>�V�e_#�jG��(�L�������?�����6Y�����{��}0���0b@G�vC���V�;��8���b����ak���w`�A�Z�<U����st�YG���h���`�{�����}뷈ɢWn)V�=ۢ��ܧl�N��F<j�z�J/�"���(���������6�+���h��L港�T~l�:m�O���%�K3A~e��UM���K�iO��������N&���G�����ӹ	f�)xm��Y���zv��6̵��e��+����)�r�7��}]F�����v׷,�0���VEʭ�	y8��u̯�E��7q��� ��K�>B�|����:&V��ac ��o�&�	_��r2�d	�z�$��r�?������䀡��S6�����/�)Z	��&� �_�����lFA'(�z^_Cr��;N�R��0ş�5�&�s��>�ؿ>��	[��a����t-�7�~G\�Ї_��(S����j���q�B��h�ܧm�1�U�p���3@��_��,����r��3S ���!
��3�M*�X�.'� l� �&,� �]���Ys@7/�8U�CW�(�1s�D�jߺ�ٷEl��*�\,��;���~2��W疣�p�[��7�B�Lsj_��S�ַ�El��u�gi$kG���B��֟e���l�ҡڴ�7}�
��?�F��6?�/�}�A�O�%Sd�c�5]�4�@7D�_ʸ9)�><���iZ��]`�
b�E���R@Iˈ`�B''���DJ8�l��3��5
q�?x'��X��20	N�!~~�}��𖠄���mP�v�t}J��(����Azp���FF�L���ȕ۔���];H�Q���Q��-g�1�xO;Rai���$�iFR���S�q�Y^@i�@-�%���}a�]���zj�� Uwj�<a�����1�g�^Oc��)9�Ê�6����������V�j��y��ǰY�[L��X!�:����T��������(�F�F��%a���h]��b��P���$܊����6�ύ��l�`yۼ�Vr6��]V7���`�bw}Q�5hX�xf
٧��>��֒��8�O��pŽ�7|X�e5hHpAj:�����H�d��7-��?������[46�Y+��d�JW[��b�T%� ��yqy�H��g"���y���٨몯w�{&�`(:��-N<��tPy��dَ��b�п;��P��E`��X����8�w5���A�$H�-�23=}�0�o��w<m�F'��Zkl��UGe_�ú���ݝ�iEw�=FZ�=�C-�8���#�Y�)1�[�b� 4��}�cy��?z���f���xc >Gi�5�#�7��=� iP�i��<Ox��K�_[���9���c*�%;�Y<J�EƷ�?gjqw��s�"��<��d��x��iॲ�;d�(�f�R(K��l�h��k0`sj�Zi����(����7���
<;�Ti�&�bF#��Lr�Iq�����&m)̆)}U�?m�C�����J��[i�yx!�m�7�^��'H����깶LQ�?EA�=�Fn�ێ�b�S�ߝ�:z<�)f���lX4��τi����.�ע�$%j$�*�?�nX.9gh�7$?u�ع��՝!5����֐���`2i8�k�ҷ�+�5t';X,	�z�&� F���F���
��L�E���[�b�����X'>��q���ts�؇]�'�?'D��/\X�8"��;?����2� ��Ft��g/�m�|mC�t�j������Q������T��Ճ�}u�����e��	P?� bh@��A�=�f���|�b5�����B�˫�0t)�̉ 4ϊcz1��׾�4�
z�X����X,Z�e|Mqi#S=ED�&�UbɊm��rʟ����X�^���O~M���X���i�J2�����(�2*4�y��0G#�F�>R*������\u~r^ቼ��%ǟþ����a�����I{@3����O!��З�^)tÞZ�ҳ�5Lt3��_3�P�Fz�z^����іfBP��kgA�2�8O�5v�MT�;����
#�NU��$H%@�
ޫ߫V	5��l���u4��"�;�Oԉ�S�+em;�~� ;zM\=A���d"G��q�Ӻ�b*j�{^�����6p �����h�	3����~�v<��뎆`����#]ȵX3%Q �v$I�1��	����.��f1r��o�,��P��EƤ��C*���'��Xb��;����l^½~���=?@��d�J�K�uë�3#Dj%N�_��3@у�D���5��샩��� 4t��S;A��N�f��9�]֟<,ɼĩ���iַH����_��:�*��O��v���Z��=��� ]���'�)+�9aZn��Ʉ�{d�8L�)v+�<ݯ���?ڎ�$�n�^�N���X�����4���6����	�h��9�&g#"�� f�9E!�i-Q�+�e,�T�L� �T)"�ܟI%"��mF�X%�b��,ݽ���Ǣ���2L�mܖ̳휳���f���lE�7.G�϶N)��L�|�
���	���PSy��h��W�k~��e:��ad�+1+9v�So<��4��8��YW�)�oW�ɚ�x�'N0�I��T��s�{[й�Ov*���v�����]졻aφl�����g�jp�|�i,^�E�5K]���,c-ÎN���iqxƒ1��A���9t�h�y>�B��KF9F�[��Hگ*i�h1c�߃��Y:+�E}�O\��A^F�H�C�恲��J_e/z|��lL��*㍌��P�?��~����\F�8���!��J�߿� ��όv5�	'������J�^�!��ac�Zۂ��]��GM�:�e���p2���ꗒ?��pܝ����&������(�u9��H88]�ҏ&ws>����;����~�v�2�c�����M@uc��)x8��&�?lb�� t��JB贽�@�eB}J��s0�1}kn�l��}���@����g;O��SR�Z�_r��ũg�����D�I�Z�e)�Z�T�Q6S�J��Db�
�=Ö@c�}RZ��1�)#e��G�yl�G��dQ
���v*�"'�`=´�7�$%��5�:B�14ݻ7���4���"Xd,�k9�}�� ������f|`\÷��zx��Bh�,씤#�(z�>�Η��쐅��hcގ�lq�$��3�A��{b�hJ����f"WJ�L�eK�W{�iz~d�@i�n']I���xJe�O�X�f�&�bo��eه���Hs��0�B^��D��^"�]�X�"羪aC0��K�5���nT���Ju�l��c��[��h����Đ<���6�♭�A���r�ɾ:j|�f���AV�˼��3��iv�xp���f�bM�6Q0�&>�����E1SOH��e���h��g�Q��A��tM�����4�#���oXlxVHYEB    fa00    1950�!���ĉ�L� �E#�}������ЎW�3��R�9�5 5n4�wb�-_�2@~�;ę�n<D�}w��a-��/��A`�]��l4T�p�M[c%��� 禗`!�=CT}xB������^��vm��E<r���T�T�hfΔ�stJ�EI9�V}Z���T�F��E���=�NI	eٸ�_k��?/��p߶ǧ���n(�Yڶ��� �}�ɝ�>��Puâ���h�s�S�kd��KTp�_�����X��/�����RBW����suu���#�Yw5m�����'CӇ!�f%�?��:"�ّ�!�a��<����"۟��<h]Q�s��h̯&}��1ˀ��ޑ����o
 ��֡P�Ȩ ���~�D=}8�N�
��A�:D<H�s;킾f^�����.�z���j"Κ��m�����m��ddz>g��"�&�f�;Ѥ�XNm"�MMт���e部��i͟é--��ܤ�ЌXޚ%w�] �%�揋b�L�y���>la�\m�\h�I���D1o&��ꘫ���x�� @�x2����eW�p�NN���\qM����LݧJ���5�e����[�QK�VjqߵQ�M019y���"�Q��4�えE����;�A����0*�tZ�����+N6ނ��6A`=|��c]��*;�9;*"ȵ��a��XQG��df��-k�����c^���ٵ�=�����Q��RC���բ�-����]A�h*z������cG�����(�h�d곟�����LDso�d�Ȟ��h�?B��X�4��϶;�f���K�V���C7�7���(��|\�v�Ũh�Ctf@S����=U�fbRKf��@6�ꖯ� R`PM28���-�����}�)���[����C_�ͻ~��g29�M�c�X�v�^a�E���p��ׯ.�3��<�<���	h��j��yg¯�y᧒YB���W<\���Ϭ�y"2$06̤�Z����K�c�� &��Mnvޮli�0�Zپ���>��#���;�z�S"~��K�8�����`;1�+��o�9�9�FU�H뭸}�?ag5���}���L�x��9ZKgSG�ƫ��&��;�^.f8e5�)�HO7�+-�3���oG��Hٕɲ���#X�#�E���Y�H�4q�Md��x��VA�c�	4�|���iԕ:����U&06��c��W���P�xl��r4���\��юhZ�4[.n��'�ˆ�:�â��2�k���X�g(s�������5`é9�{dwF_��c�8C�������M;�<T���6M_KG1����yq�BNS_z���hد��E�s��D�h�0Or:�ـ�'�Yp�8OF�ĸ�w�57d��J��F_P����S�7��bT �Rܦ��@в��ʓ�ݮC��Vr:�N�+-�����(O���<t��xRS�1�i��ٽ W�\�#)Jda����zò*,3�cԯ����l��o	t�0����%jM�E"��Y��������΁"��	B���t�N�Iy�c�fԪ�@��SD�+���A��r0tO��s�{�&O�9ј�$��n�{L]�"�� ���2qK�,���$j7��E�o��nx�9�(�Y ���X�r�!����z��A�@SY�G�/C�l�EonDONV����(���~{�zט2�����+S�t��G:�Q��'"m��6�"�`� !au>�Y���/{�w��sd\#�'0��;��{jocM�+\L�|��$�IcwX�i�n���g8`~3|0Y�����λ�K��1�A����s��^V�}h�7,��A}_^�/Y�@��d]�W,G��&��iY�r��!%��@7�&'�E��#H(G�	�H�L��a�x�~�2�C���ΐ��N$�<g�3t���u5���d`����wvs��`\��t|�����e���U�O廬V&h��<��B�) �z�ep�o�Myno�,i�iͺS�8H�g�jΑ�r�߰��-��X�^|�{j�gBU `�|�)%����i�"�w`5�!g4���V�'�Z�_!��Rg��A��|+�6��T�1�R>�����[�k�W� �\���l(������F���I��J�6RCjx �,��B5MMo�(ٸ#V�t1�1�S5��Q$7�?ND����4M���3&��&������U �:-�Ԝ�eH@"G�=�f�}i�x-N˶_�'�/A��L"��Z7[�@aځ�!�$!��ِ�[Cy���CQ!�	���:FD}�^�_��b{���6����U�
}
O"P����RƯE�q�)��ҹ����� ��Fg���m�=!<�⸲d�ێ�=ϟ�L�ڈw% ϔt!�6V��׈&�o��U��)�y�Ȏ��"+��iG6U�"�ukqx�%@!���`�͋B>��{2��p�k����y���AD�z�5/_�Q7�1�t��wmǵ��_�!TPm�v+���-#Ra?� ���@�	<|xu�l�9���x:EZWć�I5��q��`�$�^����A��g,��-��g�(�<;��6$L};�2��T�YD�<�A���2�k!��,+���V	}*���&��
}�P6`����hv��Už��'VƠ�DFt��snCV"Wk���U���?�,�=��^��9靈`P�^�3�"n�:T<�x퇒���(����f�)f�D)��>t��U���w9[�>R��x�iD�F�s���)���N���7f"?� �KP~�S1b�啘�K+�ߕ`s2�����	F��ˠ5�Я��7������uH���u2��d�L��*��.�/b��:�{+3gya7�9�p6�����̭��'����0�]�l$�{)�/|�����τ�9 ��	�4`����(+ TN%'�&��Ĥ*�6i9��V[�eCk�n����O�tTX�񆥢�Ux���>��l�\ӯw#U��N+�? }�z�9ċ�_�c�'��e:b�%O85�
vp��Mh]�
,�nH\���~�Ji��H �c�+�\Д�R!2bA���]e-�pE���ڢ� �J���7&�/J��-�nl{��=��W�3S\=?F��8Nv0%8�坪WI���c3�����ɜ������svÝ���t�y���cb��_�2� P��UA��=�$��|z�b3�����ˬ�����`�y�Ȳ@<&�!XX�9
��b :Ω�����������7p�o^���`�aAB�����_�����[[˱�q��sV�2l���Yl��&��(���,x�P.R2�ne�ᎌ��z@��,�m.�a�Mտ������L��3^4T�{9�h��<�*�4����VL���!�RvӳR�^^��1#���6�$)�c��\����;kny;��{��p)b"�fw���9���s~����[P��O�Uj�w�<>���1٫�^l�O�"��҇��s�ؕ��
�X1��V�:�\o��]>�"��E��`����L��+��#e�_eq+ȳ�x���l�~��X�vg����ɵU�6{$%��V�p� μ�Đ���-B)Ȼn~>���P�+�[7R����(�����H6�yk�=z^�#`�{U�c�_4[2z�xه��� �?dg�ܱA3�$��� ��$�U:�j��uH� p� v�������$��,���
�ъDmA����6����Kn/+1{#�RQoyo(/ܢf�DH�#�䭀;�x.=y�'�՝�,B� U��R��&Z~�<ӇO��w�Y�H��T�:�>�Ƈ�u�{�Z�6�3�D-k �&+`Cr"Vu�1G9���sN,�F����W�RW؁��a��)��0�92lO� �c�Q3q	��\m�u0�;��I��O�0���f��V�����:�̺�u�RDe�{�fhV�
=p�TݓNYr��	���0�Dm6�Ei��@�s�V��	]~�&C��~�ｦ	%�rQ#ہ|6�c��B�|���OFu�x�H���:w����gRհ�2[+r5-y�3n���.��9��9�\�'��^���Ъ���g"(t�/J��y�\5C��!QctUe�7�r�r���:1�6���\L�;�Kv��x���]F�<�Av��]~Ш`"n�<�q~�Ѓ����8�9j�/f�	���'ƅ��V�8J�e��h�y� �`����1{EP���a�.ƨ���R��h-���'�2DP)���X�4`�I�m��Z��K�?	��yBڜֱg�b	���<>bk���)-���=GOD�JF�ÐP���`�����G]��Nt��?�/���CH��~�����䙑��Ѷ����(��4y��k=2ˍ<��c���)_��{	S���_!6�.��a�c��$��� �c<�]:kLDL�������Z�E��[�c�T�u�d
���L����?]Q�n�N�w,�_#�W8��5�\��?F�:]�PޱX�����,�N�pe��Px�J�&n&S�C��^S��6��4��Z���$�I�E����l�����V#��ӘJcJ�4w�{�9i�E�3�*h�4���A���+��o�RnR&<b�"�Z˅qf�
Vu�h%�.�]ȩ�e7EM��'kO]�.��|ޭ[��]���@Ƿ� ��)
��{�~hQ�q�#���=b�g����y�l��j_+=ImO ����v=K��$������@	��T��{���k���gDK]��EsI.*K�� ��L(��E)�/���?�F���-�����?6[�����`ǣ�!ɭ� � ��u�!T�*Q��&?���6$�Û�KKYz	<��(s &EsS����$>�X�<�m�	A,IB%�t����)�Q���~���u�aEL>q���j� ��@R�Ф����2>o���JVGך���!��ap��N�
���J+�X�wh^�`�A�!Pō.�l�Y�9�ף��"��yd�x��.�T�Y�����"ދ��o�^�ӿ�=�ϴ�E3���-��^U�����{�d�ء
(P̯ع�{ �{�kv꾸O��	�n��O‒^�w�����13��^1O�.g��ܸI.�%�_�ΦQ����۫�w1t�P��2���f�%�87(�]�qX��yL+��w
 &%��0����IW<>�'�#���)�_����O���΄�\QC~²��ڃ2� ����q}��Z�ޥ���/X ,'�]��3rj���N��
o�r�:?�|�ğr�@�i�p�F�&*�[zX�C7_�C�&9ʼ�Y�Yp��DF.� 3.Z���1���������l�<בL�����.���['s6���*���e�?�"W�12z�E��Ɋ������W?c�U���Z߳I�'��z��������/�O��u�ε���Wa������X_�Ȧ�>wn����o��/UQ��*�,�,'�824�a��Rz�gAEF�l˽��<����Q�Kz�n[��|\�xY�b�`�qVE�K���htS���k?��E�Lp��"g�~R�N�>��;��O������qx�I���ysi�"L�p�tRQ�	1� ��������,Dq:)8�R���Ҽš9Z)����_xv��k`��j��qE�|��L�{����7q�>�^����LnI$7�bm%�Y*�e�;l���+�����J�R
�9i�K\���rKnllzQ�љ_\y�V�_��j�?>��9���h�a�={���
�_{��rnP�D	���V˽��y</��F�]w�8I�_���}[��6ܽ���`���3�Ӡ�N3/��8u��-C]"MX��L�P�(�N��P���/U!-}�s���O�"W|)8�mStꪧ���0�0��I ��įb[����вBX�p�M�����a��c�C -��&����8\�q$_<v���k�4����UI���-�խ��-����8�e3��栖&6k.�MYq��2��Z�wpHP��^\�|��-���>�G�c ����
\U�&�m�5�eF�R!��J�*Lƻ����<Ԕ�(e��]D�4좞��W>���H����N b�C�|��w�����j����ڝ�*ɐiKA8�a� GA$@��-�ˮE����S5�;j�P-����@ Ş]�2��7
�����=�+�ۚ���jbe��N�L�>&��u{1Ԑ� �|��m�G��T0� �������ΖH*�,�Xm@�i�]��u�����(j�ыr�
�C+ܪ+���p�����͹
7K�ܣ������e��Y�'58��Q�[%���C*]$}��-�qrO���Qڬ��HC�_�w��-,�@c9�����j�����UXlxVHYEB     fa1     440�4.����������8�C�_��bK����q�� ]Oȋ��E��%��p%RDC�1T9�if��S=���	�3cߔu�o��|���ŲG;V�,qEQ��B�hY��O�.nL�� �����L9�MP����B4֜����
q.��z
�!@>5{i�D~gf��m�.�s2�-UGY�J�~g�F�b}s�Xw:�į�A��V%ik��|3x*�lK~ ��G)��-�ڡ97�E@׫c���eO��6ͽ�J�,R�AY��;���e��@���y�[%s� �A��f�����%�^K"t�����M�!��J��J�^��*'�4����h��&��v#�$�a54Ilgm���r�}��%���׏�"ȐD�����d����spyÃv䓄�8�|ʚ������G[��l�ڇ���0�]���g��B;�(j���,�d���Wt6�$o���nћ=�
 ���yw��`��9wH���J
��С���M[^MF+#瓸>����+2�s�_�E<�q��2����ښ�f����y�B� #7����)1+��HH5W���
g�w��$����D$�RJ����ܔ"Ph�{3���>��F�f��
y��$�|x�T'v�Uw�A�6�̺	6�$����e����A��3��ھm�p��T�E��ֿ>��O��hL.O%��L$1��$v��Ez��sejΌ$M�� �I��D��g7vm�_K�s[�z/gu�g*�����^'���gU��:�c�rs@��P��Z�-p�e����L���y�BG�WB��ae,���قn�{�r��~sK�������m��7�W&����Nև.�}DB9 ��_.7���h"��,��֗��sѲ�{ɦb��x]u ",��Ō���L�ZH*���v�۸l˞�6�)����������	 ����paD[A��aْ�$�_
Y��@�8��!}�w��`g�'�"��͆O�)F8�D�hl䌮�U����4ʩ���_ų^�!���p���A\�l����3�$��bq�6�^;��	t�S�Y*	;\g)73�y�h��`�{�.F(�1�G0V�