XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����H��毝����O��s[@�e�X�þ���7%I��A娭+\�2���;;�D�aG��Y9��ä��[M�Ќ�{�`T���Eq�Z9�VN�h:��7���a��;p��gP7�+GV��2�x���o=�M��˗�����e8�C� P˂f�!�/_���H���>a"�	{���T�]x�?ZG6�*m�/WW� �%n���\5�ыjD��_��E�[A8����+d�(�����sg��iA��˵���塐� H��������|�}PLf>_)��.�q�/ μ�Y�KQ{��r	٫0)e�e�y���>i�ٱ���r�w8<f�4+U]�8�߲��@�d�}��6�G>�t�S󽟡hMO��K"�r��*T�E���Y�p����N���������G���[u�m8�8�E�Н.�R���
���e=�m(�L1�TZ�6��p 2�.�g^����8����Oe�p���}���҃�@����X:e� �$s�tlm�6{�0�sM�(��^�U�p>9�ٸr�r�G�� �n�*�������~��v?�K���-gj�*���J��R�1N��FMk3�� a ��H���O��RKA�ࡓÕ�R��1f�3QſщN��	��X�3U��P�T�X���� [�`�Ü��s7]\��}|E�+�;Zsz�f��%�p�7TW�A|�G���k�y�;E�IP̣}�i;��J56�
բh�ʽ�fq)���yъ���a(��ɉr�fXlxVHYEB    991b    1e70T�Lj��W8�L� o�7Q�"��˘��2D_�W��R�ci�Z*]�Ջ cU]�N]�3,�1>����M�5�Kٞ�Qh'K,���de�}�6az&W�mz���n�"BT����kjQ������#�\��!'9w�����T�gkG�[��{�����A�2̋�*&�{�
�{̩�\|�C\��I�M<G��'�7`�Q�n'!�.i�y�-�g�i+d?��u,g	i��)oy�JA��ö��Z�b٣����^��d�-!}j���T��el�6�>'[b��g��<�$��H��mGX/��%��K0E�V"[2U�n��N�J��D�_��-Gɓ��UK���l��\r߇� �����q��ɝ���)2���dl����
�L��*F�-�7]$R��[9�u������C��@q���?\�;��Q��j�|F0PM+�!�x����k.�z�W�rm~h~�̗�"۞���,��늈1W���9�!���7���T�<k���$;��t�s[���숪r�����@�i)p���C�Ι޸Mژ�g����j/&�R�,�4k��K ���7N�VDԕu����+~{�'�  �����1�?"? �rZ�� ս(�s�HB������c�2g��GzP^�0_�"��^�b?�S�q_�Cx$���;G�G���v�\Ĉ&�x�)ί�z[��?����쪼�a��mM�rKa7�M
����d��A�f��+���`o2�}*�Dh��7���s	��/��2e�T5X��9�'@�&���ϩl���S��m��ԗr����bw�����S`��BE�[��z������%�hd�c�o�2 ��2���	H�OF�%m
�!�7PE` [��{I
~��7�@�U�WƭSa�����zu����a-|�.��J�~��A<4�Bm8&_�Z��|�?�r. WqYkp���Rb�[��VuY���:9��ƾ?ji:/�W�`)���́?,'g%MŐJ�`�����g5+�н��q�@���Q	��5:�)I����F��4�4���Z��!��o�T�@,��R��m�w��iDQ��7�/�:�f�oem-�"���-�}v4����?��-c^y�8���2�-�B�wO	,˘p$�d�\D1~�0L�����qZ����SQ8Ѡ� �c���CI�v��e�|���	�S���$YNw�@�;�u��S��Vf�#=��6�>tU�������C�A�#���i;���.ɇV��NR���]�s���u-*�s��x���|������
���(@�f&�2#� ��;ε4���>
��"�ҩ�R]^�b�"��݌�K�]�
><',Ȫp�iw�y-等�����c�.�:��w�_�j�࿯$�VQ�r���Zv�,c�+�R�BK@VZ�4b�Y��G��'~bl�����|�rUA���r����t��m��v��.*"���$٨���	vZ	�^�6pp�:^c2t�Y/���BK�31�;�n'e������+ͽKθ3�̉��fפd�����]5�ZI8�!��;L��.:D�!qvD5�X㸒y���=x�M�OY@v�X~:&/k>�����	�����fln�'%���8�z���:����fFq���2(����9|����o�i5�tlAenhz%�e��DV$5���$<Zn��C`�$�"	��4 y�)�`l�a_��1���q8r̘f�0�L�˿G�X{��� ?�o�Gr΂���������9_�]�J�zz�y}���J(��=��J�A���w��v����R��bv�wդ%i�E��x��w��m�`���/�)��b�
t�{s�u��D��Fq�sl����PB�\¹�K���=(Vpd��˙�����U�Kz�$��?([n���\�}�v�q�&���BcH��KgB\=(�B}�#e�{�)Pu�q`��[�S�w��Yݞƽ�eH�κM5�6�����g�� �O�[�ʟ�}�3��˗�J���E&@g�!��ZY4p���n�H:%��cR�G ��M��O�4�����l^y>i��ff�ۉ����v.d���N��[g��45��)���-BԾ*Ym,�'��3�������n�>�4��m������a� ���C7��s�)�fw�08��B^�����h�≈�9��h:^�_ɰ�>�<��̻~�v���bDG����D��Ҩ��jJ+�T9�h�q%: �Ԯ�p./�=�dF!a�`|'��&Q˞������l���VJa��O�i�C��\��/�zg
�!e�P�G��|fh}�K���?V��&·k�ϭ��W�}� ��rw�)�υ��3���v�7��,ء���_�3b%J���R���Uf��ٷa�耕�x7����:v��9-�FS��F&�1�����˞�&����� ��yL��U>l?��{��!ċcFBv:JpQ|�@�}��'0���p�SI��`����9	�)�}�W�b�^K�!��� ����a�J��uK�y�ɢ�{�ؑ����.+L#i:��{e��n�-�Q��������G	��߽����Exն�6�+�Bh��*��-��9F�{���4-1�p9�˙wb_u*qSS��@�$�AH)��Γ�i��ˤ�4���6�������HuF0y�}!ȭ��,T7�to>�vޱ���LK/.������vu��t�AK��)Τ� V㈭R�v�b�$���fj�0���t1����|��{����6"G|� �!�ID �-�
c��h.��/N�)=VӾ��u��O]�`L��5�t��C�I�����V邈��r���p�B�x��6Am@xkҾ]_��;��ȵ�+7U�ymbۥg'̕����6NEHR��
cRc�:�Z��Y���}?��S��=��R�6��w�m7�Ry[��20M��Zt��LϨ��_\��1R	ںsM�;�Q��������©�rL�?@p��hg�hV� 7�1g���"��v�X�F\�=�B�o�"l�N�"�N���dX�x���v^���7���o�'����|N��h.��Yi��ub��`�w���x	���㞢����:�������/�@P�IM�}w��D�ܛ��Ks{�-��kU���������s���
Җ��纏' yr~j�Mх�@@g�d�v����?=�+;)�qL��"(�p�\v��]\a�@�h��� l���m\�Nx���0�?�!lvԪ#4�e�*��-V�-I!��Z��1�zM���թr���a�����X�	��� Q8��6�:.>��Q���Ӫcx+�I�%&���W���.ˬ��-����3�
p�-��b�U��)׈�����V�~7Z��pbJ���� r�V�ȫ����i���%`��f�I;U���Ȕ{i�O��oWn��}uX���d� ��c��H~�2�ͤ3o;M��s�H�k������
 ~u��RF�L!&H-�a	s*�b�;���� ��j���\J�O� '# ��#hklP�#��Q�����+9���Ρ�B��6f=+�v�{���y�����u���FE^�3%Z����ڵϜTae0��E|�,�i�o���;T��{h_�&Y�8�����5��	]7Y{@����2���������}T�^Ux�Dޘ��a,Z��m�8!ҹ]:�+��܎�T�;`nqpQ+S_����ys���H�<E^�IH��K��_�NO��6��0�j���&���lJ有GK��d�ҳ�h ��f&	IUC&u��e��!�`�K�n�-��q���ϡ��wX�������i�V���K����ː�SOu��ڲ�;���U��A<���O�fӗB�FMCF��l"�����^�P���I�3���bs%W-�`�Sk��ޔH�588{ˈǗ��$�_:��:OQ���_$��G.���S��=����#��Ǚɸ��%n<ˢ���cX�,�c�i���od�D�-I��	��@ (O��{���_��-�U��: 5Ko��;O��<�B]Y�˜]� n��0L�n�˻wR�K�9��c����*��
Ue��uf�ӏ5�9u���Ζ3���sq�+�׫i�`d�PAXٶ��×"oN�L�C��B��>�U%��!,����B����mR�U�����\���n��O̖U%��c
$�����}�/���x��(���G �N?:�m�?%�˱%�Z k������m;��Jg���u���(NrX���X@���z�ȕXlcMй՞�QB�(
e\�����|�,2�	�Q��{�� ��@���]棗����̟�glw��Vs�t%8Q�+\��>m��P#x�"�|�ϭ#�{�7u�]	#����Z�@	�'%+��bA���Y^����<@��%��
^���X�H'X�>>�"��^�w�i�񜲔g�:��-���,���s,r��̡Ah�ZXx*��fަ2�(%cK{�eM/`h�KJQ�4{�nF��@��G�a�%�]���%Bc�¡��5&��"I���Y�Ey����V���<V7K�w�1ǳ�uyK���}��Ebl։�$`�^�-v��7-JĤ��w���m���Z��Saz��ǣ9�aChX�=����~� �&B�7�P}
�r3�tO�J8�}�r���1��6�AE�w�P������b��׬yx&L.�w��%�ʴl��ơb�{+4�Dd������ZR|�f�6�i�-
�rg	|fr���z�~��m�zN��ۧЭ2:�yD:ڳɒ��9^)�k��|�{l�2���;��է�Ƙ���܍��C��&�K�$� ��L��aD�#�(t��A33*��"�ı��eIΓ���6Y�)�ø��6�=�
�RސI��8����.�c���b.��؃TIl�KO�\hV���_v���J�аF ���|f�=W�jԮ:�%O�О�Qо�C�H��������U��A�^k�X>�[�A��#��F[��5@E�� 	��A�(�vH}?����|�,j��W]�y��rEO�VXp9�[��=�`}��&��3�k���1Mh����[�*wD��z�{�.� y��w�	xaA}G���@K��Y{�GzѢL����Cv����b0
?;	��X?����d��)}fA!؅$��IthvM�f6�ЫT�ݏv�׼�`��Y��8�D�$K�� �m�)Q�Bam1>��`<�m2��i8��12��<��$�5��"�)G0L2+�a�2�!�.�.�M]�Ӑ�P�J<s�
�Vv�L��HՅ�!DBVJ�y�+k]�V0?^j��{"�r�K��D����� B�'��v�O9�B����"�u,b�fHo� AK�U#9�q/T�7:��n��@�1�X��f�Mǀ B�'jt��4�:��N�?��;]���a$<i��	�m��v�1�ț"�		p�Bq\�D���������K��ys7Em��*�JL,,A5������M~�s_r��_���z�+DXx{���!�V�1���zS�tj��3��?�۸R��W�����O2_�M���x����qO�������y�Ӆ%�(��ܲ:�K��|��������M~�{M%��V�7�!7�u:- ��47�ueJ�/���
z�]����Z��Dvd�QJ)��a>K1��s;�/�ɾ5z>� 0+�@�x���=`�˸�t~?>�]��㔆y�ZV�����\��x��$o����gx_#��	���f�b=U2��������Ƭ��e#��Ůً Q�Ԍ�H���q���n�BIOɀ` 2I����?b8�����S�YGkm�چ�Ϣ�T��i���&��pq�B֘!�*n�G�$r)���FZ��P�ۄ��ź`B���ī�@��@+i��@�����v��͗��H��-��vphOӢ5E�hUf ��+�{Z�Я�5dգC��'\�x��m�Y|U�J�U-EWJf����\��>x�e	��"��Et�e��ӫ1���𙴓����*#)Պ�οw �]�#�g�u��	=�'�}ہ�h:�T�jX����{�Q�'�M�:�R�0p�hUY{59���U��l��p��~q�Z�FU.:�C6{��$/��v��x6d+`0\`�����)H���l�rV;�]�*��ݾpy��i�o����}m��U�~�V{�[�6�N�?f;bWc#��xRٻ���>�����>ag>񤽜Dc��>�l$�
��5���3�x��0ˆ����%1��jM��]��y��߼�#=L��
F�G�����{�Bͥ�R�n`#^h{Q�|�L��t�L�gH��ia�`g��E�4�pˎ7{��v�Jţe�ŗ��wÕ�Sյ�Qh�iM#g�cjr2[D(}�D���|>u�g�N`v��T!%��JT<�"eub#O�qm̸�&�Mɍ��'�o
��Tn�CZ�)f�v�;���g��5ʻηm���3V�C/[DY����[^�(M�9�T9�����:�Ǩ��̲�Ğ�L���-əJ�,��^�!3;��E��3��<9K����c���\�WY���XF�Vs}�et�<�-�S4�y1L��`�Pʷ�C�I��su�ݬrLC<��g1�2���ET�y᭿�
N���,f�u���!�Ԥ�[�gYv�tn�
=_�\x��Cܾaja���� �x[�����M�toV|t���9:�jk���N���dE�L��u,a��ä�2$0���c{�KjF-i�%Aɏ�I驭���C6��:r9H��Q��?j�+  F��Z_&��+bi�g���ѵ�΁�MPvչ�+0햆U�ö��Z+��fn��N܉�^ *�u���~�RC�1���Gw����>�rɋԚ���km��H����ӯ*����d�����"�i����C;3���:���W���+qh�M~�EQ�U�V�I)"9!^}"<)�x�7�d�}>�̂�W>%��h݆�azb�L%�.�L�s��f�Ӯj_Ғ�z/��|�� ��,b︚-}Q��.��� �XဳU�$9�Pdˣ�M�K��CF	��Al��� +�6���z�2IZ�4��V���1�A�N��"�0�֋Ϥ�M{�&��J�w�a�o�ڰ�i[�J��\B���,�~�[�\�%�X�Lo�GP���i�.�ױM=>H��M�A�A�v画�59L��"��?DM��qd�	| W0�!q�����/Z�� �u{�[J+�p�3.�wϞC@|NN-KP���~)ᢡ������h������<̣<��=�e$�Ž�����q�Vk��lV�
Զe���[�4FX�El#>p� ��#@�M�]��$�+��u;o�!q�W�\)�|�F�M�Iyg{"~5L�Uc�.h�1��cj�s�L�sV4"�>kB��/�Vg\}�xf�|�iz�z,R�n����Wh�#�
�A=���W	(Wc;�[� �`�h�T��")�t�V���,^ 9߸w��*4$Ё���Q�����zԆ��U�9F�i��R�7�j_趐:���O��1?F�O��Z�?��=�d��jE����b�a���_/ơ�_��!�ǔ���%}rР��6!7�K��IOW