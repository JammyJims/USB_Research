XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bW|���R��o9}\Yt��"NP��p�;�e�,��N��!��ճ����hM�i�q��^j�$��:��+�B}}hE!�IDC3g���Rrn�\$VdPu	u��)np���G2����RSռ�iט�t!��F���$R	*	�iv8&�(�B�;�e�*���6ť���Q�gF]#�ϯ� ��<6����s��e#��+�R��)&�^`��h>�Ep��,{�}z�	�ѹS��$83E���yY9����ԗ(�/������m �-�;���%�R������i� Y�re9�#8`�8��������(A9��Fb�'���e���-��8Za�`pc�J��%�T%WW�Y8�G�6'>�99|��q)���n�v<a�lv[B]�{���4����$�����G��A�����IcHI�@���M4f9K���%�5I]>r�9���x��ee^�ȼu7�i��5�2X�b�4xRfo\�q�(��A0�Q��R:����{;��(9h���9{���7i\�B¹ 32׈���=4y�j�n�W̶FCӮ�������r>���3�k��%���6L#�a}}�,ʚ �������{�l��̑�~y��+	�]R�(����2z��NҼ���.�½j�!���4�є�k�V'�K�~��0�	���w��3T�Wǰ~[lΠ�-Z��QP�0�	f�ꚭE��hTe A�9]<[Ǌv� �����Lz��U�����g���I���I��N�+�����XlxVHYEB    5421    1070m8o�)�� n����H,���(�i��¹г�=������V	��p0ca_zL8T����{��{�2?V��h%�/�H�=7!n  :��̸�
�JԌ�';p�~ӈ-�/�IPp�/[͂%�SF����t^u�W��)L�Ұ��{�ߒ�'Ħ�~�:���L��.�oO^tagJ\3\te=�O	T��ܻ� ��y�u֍��~%~%�ց�������h��LH�9�<�����|��[�ۑ� )OK:�����䨭yR@��)W���D]��(2m
����b���FT���(?�n6�@���>�����6]C��V������6����H�I���Ie\S}9�nJK�j����sp5 ����|�=�?$a.i�b}6��r׊J�[B)f�!��~"wT>�;M�7��]��ґ[��'���u��7q���Q�3v�1B3��;F-�0Xߤ����*t�Du�l���tk��ϭZY�л�h�ȹ��x0 _Y�s�O�����ǨW'��$�/!Rg-���w�K�&�����I�`���e�C���Q�oxv�$�8@Slʲ���s������S�-��7�bɡ�

Wz����c�ܚRԳ�K�l��Q�]�0fQ!	G�h?�F��Q�C�������)]?�J�c��J�P;�N�f(@���!
��3����#r�cN ����%D����H�o
<���n��Ѣ�{jQ��|���XE0Ֆ��ց�4��`9uO�xf}lw�|Tf�*��vG�í��ps��G�C�P��pa�B����=�Ћ����ȋ��!���?��=D�$;��U�ѷh��j?�F�n5��D���}�lAD|,+�����İ�YJO��}%�4��[�1��;�������4�GXKA�ٰQl��XkA�:q�H<,�]C����������`@����.S�Z��a�JZ�:��̎��?2��1�؁K 猡�]����{���X:�^�Y&�vSUܓ���W��)t�\ɢ� ��]��4%�'�&O>`�hL�ޥT��������E��)�B샑��&�ݦ���4�:��H��,�O�*bs2w��r�j�=�}���w�rk\%|�3AF^����9��N�mY=�٣�F�Z6������	ڌsr���"T����s�פ���9a�;�菳��E��w>2V3��뵅 ��i��E�,� {��j��=�$�̂׺�hp\ho��p_Bջ�#�(0����	��)-�$ߑ.�C0)D���`#ghP�L�+]_��5*�7�m��Y�4H#_~�y����6�؜�Z]����´����e�v<(�,�x6:|!��Nȃ��n�e�3BD/ ��?$�N��Bak��+P{a��ܾH�$M������	7��g"������(��d�@� :x�
���c{ĺ?Z�n9��5�91b+���b)+dB���VX��_�ŕ�~�`$MH��W�X�j0��4��k���̡�^��~pc�������hx��qXt����� �󞭖_ޖ��]/u�#��խrT��Y6i�*�[��X�	H����l���T�.@�A�y��A�ᦔ��%�ײ�X�,k�	gI�Im�
�vlh|����*��� =�(�!���ћn����ڱ@���"�Q�y�y� ��1.��b��6X^	=�vuۃ�;�A���C����5" �4ˤ�^�Xϩ]�S��>�8�י�	�������BZ����e�ոzX,ׄO4��B�Uv"�ނI������ ��l1�V'+˙q���t��$L< �X��⢼�Om��i�]\�4�}���\4���L�h���T���2y�p�ڹT��[����p�EY6�(�c����u�؂=
"mg�>�֍%���=\3������W		�iW�N���p��M�0��Vo�P��NMdT�@�/x�6�Bb����C��A�DdOD��M���&�g@ؘ*Ш8L���-�̸�Qk�~��q��+Se?�[�]mC�LC'C����}��PBM����D�Fɳ�Li���*9�J"a�k6��S;�w^1�����n���� HH����-w��w�rn89fӀn�j��\����i�m�5&����>���"��O�be(�Ҕ��A�f��)n�\"|�58��B��V�|\�5%p��2>t�h|�x$��e��`�C
�QP��B�L���C �V�fEF@캴˘���8bM:�>ӆK��a@Pص�+���WS$���e�9�+^gHY�(��k����L*�B9��nCl�m>�A2��W���ˎ1��(�\�qXc� t?�SF�س��.������k�)�k"��u�}�j��<kg�����I��E뗉�>�T�	d^A��6����=��%w��
�:d%x�v�x�}s�>�T�,x_#�c�k=���/L�|�(���?��^�����9�R���b��.�a]u)=�k`@RV\�$�����������NX��><�z�w��r:Ԁ+��g�#��}>W�� C�m����f�����[�I�b�jd`&�'�E_)��ٲ���g�Z'\~��5����(L�z�3��#�	?�z�t��rŨd�������Lr�47MH�-�A�%BвP,��tT�FX��M������n��H�5y����I%�1��r+�]V=��p��{���^I6ϳ��a=5mP�g��b¦T���|*��9����7HP��)0c�y�B��㆕��A�b�����U䮋�i��h8�R�xlh����A�'�C���__yx`��9���nT���^�7�FC3$�U4���
NR%(6'���� :!1�L�*bk�퐠�5{���D��L��P���߆)J��;��W��k�����k*�Ҡ�T9�.+d���6����"�Gl'ؖ��8����F�P8�x׏��t�����1|�Q����5_5,#�mrVu=r4Rcu�>(3T�p>��\��(��&;�a6y_�T�z�;d!qB���˙Q�-���"Ɨ1�}�o�B�N[k��;�)R�K�/ƽ���F1ߑ@�s6|���p���1m�T���-��J���zU��V����}w{�q���M�d޺/��C�_������y�xߤ�B?����,j1*�� j�o;q�����V�ɣ�)�	��#�V'<6�Ƶ����Ӭ�B�]�k�wi����}s�W�t�>%;��;�}��@���5�i�A��	xj��N'שj3�@�8�jo4ӏ#�����)�5�kf�%x��2�=�i_��Kq$Z���W�0�����G_��d T<^g�:
A�Z�5���^������_�5a��,����RaY�4הa<7ΤYGpſ�i,6�!n�i:�3�=h��3�"Qy&�g���sl"_`�S2�I�H�@�����)gH9yQ�RZ�a�d"&�r;�`���g��9�i�όS�MG���aR�h��+*S�!��4�
Ч'�U��k8�z�^o�v������j����=*-�7���j�6��$�GN�{�z�	�%��_��X��82�`a.?����_��<=ts��J��H[ �	�UZ�[�E6�K)~�>��y��c2�7z�����;��ɝ�)�J�-Ç0�sO�ަ���@�G�L ΋�U�.�v�'��u~�JnMh�N��B.y�Ӳf[H?JZ�0�W�Y�7P��f�3{�0"�&U�T��Pm�}��*�r.�:/C,��)��u�ԭ4L�
S^��ʽ��x�0FtɷN9��Y�#�����G����&��#lSG�-�{�(q���R��~va����'�<"vе�L���tVm��~�F�i�_���+ގ���	�.R'~�'�=$>"E�A7@Ѥ�ŧWĻ���| ;c��xF�*�� �w85%��GdW�9α� �'���N���ئ���Clp�u�v�a����á e)��&Ђ�,RNk�ǣx��g������1Ȉ�l�D�`q�Ȅ�q-��DE��X�߯ 2����m/Δ]���K��a'�l̈�~��eN�i���
D��wԻp�牗�^�$��p�k̦>7U�����O=�zg8�Z�ʷQ���]�