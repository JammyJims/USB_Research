XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u�w�y��;8��^��r2��5��z�����ʱ����֍0�b��Z'q�pliĄR�;��^$�B0�Yh��>�z)t�� ����]VX�ܧ������U��-��G/�Ock�VT��uL꧐�X}��X�h"��ŚMhڍT�gR����M����	p������חNZ�1X#Gt"����'����J�m�h|��3���T/�s��� A`n�w�q�)�0D���!��T���Ǹ&&��B������$�:�A������dN5sm��6m�t�xqϗ��G��u!�XB0@��x�z�N{�����r�i|�1a����d�DľuV�!��>bS��e"�S�����e��>�b \M�?8�o'��Bw{i�Z����R����D�����4�Hq�*]/���K&�A�O�]�S��f��@��
�xi��AQ��gz��ry/�j���Y;
b�t ���o�oB%�p�	���:����?g��[Y_�R��G��c��%1�D4|P��kt3p<&��0ɛ�4L^��ڻ��I�o�Y!���E���~f���X�4� }����T�ݷ\�D{3;�9�<�|DS�-��l�C�rzçU�8�q U)�C`!�~r�!����~{�u�'k�t��U�\�]%�b8�
�aǅ�K����J��WyY79W��0m�G��qʺC�Y��d��i�y����C�m&�VK+s����V���5����XlxVHYEB    2302     b80�.�����Ԯ�%j$[�$��}-өǔ�Y|ݬ'�YP!����:�6���̨C�tǃ�!��dA�噍��?��OQ��%�X�X���1�z�Z��i_��3F�pA*�V��S����i��#���a1ɔ�Pp�W}�ʇ*�@�?����F0,�/���T�-�uf�Ǜ��ՊZt�� ���bS��J7��V�@V���]\m����*O2���^�?�(�����f2"z��LZ�k2�~G�E�uJ���*��'�]��
2f֠S�*\��j��:�bi+q�g�/[��Y�	N� ����������6�q)m�
VVwf�q�F��S �Am(���7�eF���kb���,2��Ғ%�of��z�Z]�����T&�fs�V��b�]���S��)^ow�(��ZB��3�8B�j��A�A�S���n�Q��Ҹ|!D���ۈ��ሒ.Ai	�L�'B���aǱ�h2�`�Xh���"��G��}�aC��9Z��;{O��\�U�+I�h= +��Mk�]&����utj������n���b'8s�~AS=i�r�xT{!��oD^q���.���29/b�Vs^������8�N�S�@g{ʿP����r���w�`G_��x%=JN�b���7K�F�(g��y("b��O�L�:�#y/�M��l�\�x)��e�tgJ�>�p��8{U��9�/���c�+���swd) �ͩ<n���n��Ƞ���A&ԩ��
�tU��|%�Ol���U[CuҤhf�Z��l��f~t.����g�
c51X���W��!�WVfX�3G��=&���.��ۻx����(�Şd�\'X�((�����D��IL]\��kƆ��E��ͥ{�*��u��/^=8�Ҕb�W���K"&����ٷ�kԤ���NJ����__Z*HP���zH���]�TW�̙>�Nhq_5t�pC���E"�B�ScA4V��px�D7�G0b����@Z��[탼9o\0��J��*Y��X2��@���e�A�f�U<���S�F>kͩMܭa�_�UW!W�)M�:�f�J�Ol�S߷�O�˾r-^���� a�B��lclo���O�5H����tC���5nj�j��C9" �����@z7A);�铼>�0���WX\����&N��~��Mg0�<����У�lJτF�z��gzFp�e�\�� �~�K�נ��Gk*y�$��t1�Qz�L�!��xk�h~-���g7�j2�7��V�CF����7�y0c���q��7���j�k�%��W���+���.�ě���M��QzpG\=�iY��S�X��^�U|N����b�X�VL����w���x�D�,L_�������߆�B:�x�yZ�Q[�N���i��j�Uc�g������!TJ��T�ȞHP�Un<S5%��^�٘�R8`��D�N�B�ݒ���A w��Jq�+��\����e(�|_
H!"1CR�٨F���T#ä4w���3�Q���G���D˃I�? ��E�`�gz�{<kA�Q3��*��~���g���&c���6�K���� ���C��$O��6V�;���N�~�nMm�xt}�%cU�2����,.�92� t���D{K�h������8M�"���wX�_Q���66�᎚�m���<�^T��]A	�?�8K�>���LW4E� �B��-D�F�Xǌ�
JD{&�\H_�2�\�Ƴ�����d2�G�E��<��c3i���%�K��D�)�Ԇ�"���S��%>(gSm���R"��r����t���5�K��=c�|S̜���`��h9y��V{�I?�z����J�%۵|���h��X�qX�(�א�S�O�Ϸ���[!JI>kn߹�f��Fc\�||�PH%C��I9}0[�Q�p�^\��:��GGF1I��oRL~op����&s�m���rA&ͭ��L�׮ٯ@A(��n�[)��H��Shaם�|�	��tV}����c���Hc�վ:@O2�����0����yr'�k�������n�b�p8�Nr��΅qyǆY��`�8���`>H)�hD��	N0	������5l���d������#��8�p�V}3	���`g��q���"�O�mr.�q�n~O
ven��E�8J�TO^�4ѼK��b ��/c,���kW��ֈ�c��Y| �V}� �dh�k7F���s]Z7"w�����[��	'��ʟy�	�ML�/�"�~!/p�V<y�*<[�|*�<k��W��
�MGqN
�ع�a?�0g�O���l͹I�@˧���fr7����Ҭ��]����nK�f���so�}S����c�Fyy��T	^�Bz�lT=�GN�.�a9n�w�����H"�b���z�6y7���GBI�%�¨��8\陓��ף����R2D#`ܼF6.���p�=�Ĭ�����=}�-Q� ������Z�Ԅ��|�4��诐��"z������@6d��C�����a�_��LeSno���'~`/�׈9_�D%��\�?Ү	C͎�v���~	�u���LX�Fx25n���NP!�6��+�����e�x۰�i&/"�*��#{���,�B�F�wt戠�.P���b��'c�hM��4�k��kE��_�I�=?nv�;X������0@��qv�ȡ���r#�kD7p�"K�G���¾&�W���R��G`�-y����xk��IS���� �|ZG�dm��H�pqS�Ā��
���WB$�0y��������R@�q�[���|Ty�^�D���
^E��٭/��	2'�� �����k���yv2�uã�H~�?i�CG�(���P����}��