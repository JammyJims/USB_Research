XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=+{�@��I�'6 �x�:�U���t"��Zp�����7ho�4�H&qR-���B�!PM�LF@ >�J7���}�j�(�m�u�^��q'�dm�k��P
�pͿ�>i�D�� ���J���S���L2��i�DTQ�q}�'HE�\���+�W}{��|*��f���g���a����.v���x�d	J��@ �m�u)7]5k���������B,��yć��)Ӳ����}rLv�������z6ZH�gy`�"J!����1��5�qJ0�K�B�O�dWO�c&�h�h��)±]��DD_��d' 1fT�/��-��FǗ��?��s�q�&��$<��5���r�Woc�\�B��ť�)($E� �QA�S7�Ք!1!9��QJ3-)�ѳ�w_��&L�S0L�����6?yV�ᙞN�F&��QG�53z�<Ԇ��ښr�.(�?��S��2�����<�'���Qn$҈��f�Z��n��_]���i'A91S�q�0C�\�%.���d��Ơ4�ʮy�ˢ�w'N���ʤkeQ���� �t�m3���3$�6�gp�����G�87��K%�0�h�e��d�b�"_�I:H��!ˏ�B���2,g/)-�H]��J&�h?��p���R>q�\9��3��P�̸wD�u�-�D��)b�������x�[�����
�������L`N��R\t�"��4�c�?��	�=�AY��e8|^9�/˞���D쨈S��BO��#�;na�XlxVHYEB    fa00    30f0�˦�p^U^۳�X���FN�/�2�A�#F�*��~�$�z$o�ީ��}S�h~aVq}�}Z2E=*�;�9@"pQ*�ۄKG�3�Ÿ�I}�\'a0�����8�`�s@��`�#s��(I��W��YΎ�v�$Ǩ�FWFI��n����9^����n�M5 {�KV�I7���V���r�e���<05�'T:��:y�g���1ӆ�NS�B�W\Z2~ݪ:p2�R �PB�^�_�<-BQ�WˌP���t�hX�^P��ISV �8}n����dWy��NQI$�mhgc3ft-5��B����R|���mB���@�L��S���؂C-^�D�qK���]E5R���s� C�r�PG�c���DF`��+�y�����N�@K}p�y��Y&3s�*�M��3�z]�|KE�Õ�`��{ǋ�u��plE���Z�n�";������{	q��t}`��+D��'e{�ugd����M�`�����^����9΀�m5��* g��U��i3�|\�����.B4�=Iy�Uߠ�,9A�p,����f���F!�'.C{D%��I����Q�kP�b< �S-�t���0d��-�� {"p���\��R�,�ě�_�5Y��όI�^�Rj�3��Vi|b�_�6���Jw��hLT��D�����ߦ��8�M�F]��¯s��jo;�u�ٰĬ�e�d<��B��#O�}�Ԭ�v�0��:6|FBE��˛E|�������_Ւ$�K��i'A^�+~x����E�����M�#c���#�0�1a|��Y
A������[2M�����r��}�a���x��]V�l�7"[!��Ix�U��L�q��A͕�͐�r�_�^(1P�ɫ�%ϼ֔�G��'��.|��)
AH����\�@����}�����8���5����Z�$e{�4/�7�A��f<�D���
�Z/�E]�:N���oˤ�g�.�U����:8��I���1YDZ���\�I#���o�3�*��2	5�s��2�|>��o�0��ǂ)���C��r腢��%h�j<Q�1�L�*���#\��:�Y(S��ۀN��SS��1+�z\+��s���qɬ9BB臟V b�jp�\���U:�%~Dwོ]�F#X��74�d1 '8�.fC�6�	�ֿ9�rW�u��_g�h9-���6W�x�y9��Ӿ���Pr���\�q+�W�Ϲ~���y�G�?���ߺ�u��1kR0T�`��0l�%�w�f�ւ/���!��02���[��7�␅&1r^�ȿ��|- +�ʸ	[S��!���S��.�S���F���D6�^n��3_D��Ł�xl� Ⱥw���f��k.�6��ra�CI?��fJ��$?�Y�ljw9׳[����Y~	�"�@��	`yB&�F�|zw�$U��le�v��*�ء�U��n�p�So���L^�[�g^�ʽp�{�S 5�i�cY�{�x�}Z��l���]��S�����C�	3��]�/�qŕ�*�P���H��R8ԏ��dǥ2u�sϔ��fKo���~Hn�}�J.�6��G�q�,�(����+�F�f;e����o����$?�Vk��v�e��Z:JD��ӌ���C>'�k�I�{�Zf���d��%B�{�n������҅�m�W�l�.o��w���԰)>$r�7�|咡���M����
�(�"�u��y�b��7R��>R��d� ́��DVv��"�{�w��w%rb�G@,�v!|��������I�][������Ǆ��8И�}���T�(�>���x��88�:A��x9	��ղ�\�#a0���5�O]ئ��4@���tJٱ�=\X-7��#��S�ۓG��7��l0�<𥋸C�l�`�n�-��+�[&��>��1��+C�B��ɚ�q�@��"���g�Z��)������AF�]Q�=֔�i��8���:�`�_UB�����H 2(�H�N:�,��گ�u��d*I �N瞼���y,R+}��g�sAW�W����tNm�f�,�u���N���dY�V��6�g���h��&HF	�g���$!j�j������Z<���W��'=�\!TXWI�G�I:wzTy�5�-U�P�Aֵ�4���R8�-��CS�\R�d-9`	�l)zm�Q�c�8�D	�p�A�C[��0�6��i�ѧ�^�fEp��'P����<%|τ���Z78ဿԯ�d4��:���nuJ�e���QV���D��gn].>1}���T
[�D�)M��O�~h��rs��3�:P��y�?m�����{R��Ѧc�+�P(Z��R_9&i�����~k�u����f��T>מ��a�C���o����[P%$6�{���݇�=� X���W����r�&9P ����]����U�����/#LSX�ͻt4 �4�'�Iˑ�1U7�Y6�B��b(496�H�_�)�����C1�ip5���Z¤�Y:Q�d?]e6�--'?\��FM�T\-˖r����{Ѩ�8//���w>����ym/�����*�^��8� 	���u�Nd�r�#�7��֤�<�V o�:���-/��p��N�跪V�|rZ�JY~D:owt9�����v��k~w������%^Qig��x/�p��-d�P��F���qI�>��y�d�[*����^��pnq�sw�:U��|�iD��+�ýЫ8�'a	�w#����^*.Z,K���z� ��V�<o�P���%����U(���/��/}���bƲ=I܆Ś��QO�k��D$�V���0M��!�(2��ڣ��,�`4t���C@���,mҕ���*�3�i��}1V�w�&.T��U��3{j���I���t9���i.���&cĪ�[�/�hIf����N�S�"�H ��z{oN:z+�D��"�*�D��uɰ����Cw���_��h��=�ޤ�'�8������j�A��vXLz�wؘ8M_�v�s{M%W/#��*����ftJfQ����I��^m�D�r��K
�a�+��7���)ɡ| �BU��X�aU���E���=+oU�b�&�T���L�[�o<!�<���&����ܲ�I0�98� ����D���@<����^O ��j�ֶ�g��d����9t^�ߔ?'{��@X	�{�ʃJ>7rH��e���1����d'wq.3\v&O��MxV���]U��^
�tY�}�O����rA�/�#tR!���YМ��O�(&��~����ט�ǒ&��,4��]w%��a�T ���� [>�vFj %Ѥ �p��=��c`�8V\.�%�®e����5]��P�N��'�wѼOo�6�4�%�Y4>���t�1��5�'"���SCm^���/cp��x.'R<�V�_������U�`�ýg��\�0��9���W�n/�Qh�%���6<��5D�@l��W�0AJ��?q��{4�n��,M��x�$h�mǃm�����q����w��i{���d�x#
�s|�K�o�1eP+���ֈDI��@�6�JtLa�`l������ȡ�[�:�x����o�����ϡ��|���������� �97�<�zk��ӥ?~^�U����>*�c}�s7
�)�����Z�P^|x����Fl�H8��}M�v��Ō,�����|�-~�]�z⥄����X����q����1HT-I\���H�Y��kv�E�T\	�p��ch�h�-�����zYrjÈ�Yv#�p@%�AH�Σ�7��#���_� =��-�-į�5�>2�N����H���TB�msE������do��忁��m�>�>���6) Q�p�˙" �D�	���*ͤ�*���/f�H��t�{0�o��O����2*Ԑ�҂�q�T��/�1Z���6�p�x�o��O��Ll�R>K"����>�4-)/R� a.P��F�5̓��`A�$�f{��hIn�� $���;�x��,� ͗�x���0UN��!��m�xuFⵯ�y�^����[��8'<ю<�4�y���I}gԑLڥ�D�jE��穯�An��mF�?�߆E�˔����K0���o�su�˚Ɛ=��9����sD@9�"%54Չ;$z���:ݮ�T}�!�6o�P��SO����lD���^r�I��*Ϟ�\}����i��қT�m'7})��֠����ln���j6��ʼy����Thc�S��)�u�|)��7_����l�y�&m�
�U�����"��� u0ָ����g}��p$\��P}"_'�9���BKU���'ވi��!��bD����P~�n��|�`e��Y����B#o�W��Rs��|�*��R���La��t�� �C�4�X�$2˰}sfq�$�֔�V�[�L[���ړ�'��b�6�
� �ϴ�{ii�F]���dd��k��vFH�f/�%µEe-}*F+�W� �Y�ε���0ѝ�8����y�d[E^��V�f�.��t{�rp��{�'q8�K'�d�tgH.���GSj����?"��ML�^�o*�(�	d͌��Q����X2�
0�_Khȥ��s�:�8�������Ȼ�	Yh)��Q�n��r�����֒������?�֬*�+�n����t�<���}�\P��P�;�	��G:�"�Y�ɻ�mf���1��ҲU���p��_���Ѝ ���d�ƫ�i�V����%}=�8y��0G.�0|�ͣ;����3�S&M���WT-�
E��M�Ú�A�V��Ŝ,@�y��K�[:�\զ�ZnE_�M̌G��W�P�w��Ƀ2G4�LV�#8�6ѣ�v�m&tavVQL��a��!�W�3DY�=��֎�d-�:�����l�c9ļ ���.sCҒ�z�]Qks�?��w���`Z-�/4ep�q��4�������Iby2��;�c��ɺ�����9k���6>�r����:j�s�����f�g��A��M�L{��x�-����+_��^���td�ت�͓%cP=f�6�3X� �f���V⻹�X�=$rޯ8O2(@�����j����V���7�
"I�ߋ�Z�C�����;��15~K��ϸ��t�V
��3��@�::��(�P��L�e#q*8�3�a�.c� ڣ�fy�ǻ�V�O�Z���61p챃V+����������$B�'I�ݴ���:�'N�>=ڸ9s]����kmMphm��k�D����\(���y�Gm{pSсPwY�j�K
�)/Gf�e����?��L~�p#���X�����8����4�ϑ�U򃼮��mmBi��`��.e�� �_�4�l4��^�e��m	�J�M�Xґ�;85�����+$�-��ׁ��.�v�Ɵ������������+��W�,����������N�S��NL��;�2#~BO��R�v��Rf���dF������ZL�ck��,���g�|�^�������@[���=�ɒ�Vn��ծ4�GRgk����]���a/��p��Hǔ���Mw�Jپ��^�)� �fg�~�yn�30Hi9�K������΍6�Ί��!���#O��W�G�q��2�SP��X�1���y����L|s��=�.,l�W��v��Z:;Nl�凸���E?RU�<�kjN�/��e}�1�;5�����rʼ�%�q,��[a��Ŵf���ҰR�?dt/��W3��QM���Z���G��#:;�}�܀�l%��L��"H�g�1�uFk>��~	{��x8y�{�e��;m�&�-��Vî:�D��~���bO�:��aH�3��2�_�����,�������	�B��sI��<g���qF���cO9�x������Op���~dV/_�#��Q�'����N�k�JGm2`�g-?+G�ŅA
��7v�Jlsoa��GܙR��)�+R��V�����(���]��T��y��籥Ϯ[U>H��9��\��t�����}��f�r��ޟ��B`��fx���!�	�Z���7J�DH��*��u�Qqf��#�2����N�}~h��O����#J��C �����+|��I��S^�6�pXc:Їz����3&?���(�W��Y]qO�h-t(�(���7WtiM7�c��f����
��uj�2Qaw"C	��S�&I���8e����*�r)���#�k��K0�HS�P���֯�| 3����:����r[Kw
[D-�҉C��q���U�-b�n��/ˢ�kl�~麪hz�d�]�S�����]��/�P��i堽��#�g�vdl���^���{�����^�d��x&=3��p��c�ƪD����VQ|�MfX�o7�q0y���V!�Z��Y��XbVo+^qI��<u
�R�
��M��:a�&��!�
E��1��V�iҜ&i�B�.1u�7U�%g��9�c?sC�'T�r��=(�r����4Z}
�-'���M�?#�HMp�]]m��I��`�
�H�yjm�5���:���k���8Vp8���W�%@�����åA�r҉ru*���+��~�eJb���e��~ `�^��Z��3R��M��������8�6�9B�܂�E�`��V/Z��p*�^b_��h�\����8�x����s��0G�UC>?�C4�*^ӣr�GI�ɂ����I�X�(���.J7KnSJ!��X�2�n�S(���aE��&]>H�,\�?-O[����r�2��4�u�>�� ��?_d�a�FX$�2w��$��5�7}d�]O�q2N�����H)��`�2a��[�g��6�y���H�ȫX5��M(evn%�����ЄCނ���%nįH\Y�ƚ1�����=푇%8�Fo���aA��ks��1m��*�:��&v_q����8�F�o�z!�f�?���'�ޢ����]��Уu�
��P�P�����
���k��s|�"C�����၅�T���&�.��fB�r���O/=�6�N��X��M$�׀�UR���(�|�)e�m�&7�um�����k�n��s	m��¿y@̿����^<X4���NïW��k�@a}��
`���i��ݙ�$\��/��)��$��T��hw� �h�ÿo7�&A���I�}��Gm�I�
I�(c��BH_��s"��Vf6�p|ǵ���~v�*z�N?{�,fV9N�@`6�s�ގ[��]_�9.�cI������[��?�;@"�ω������_
~��:�������+����C�F��J��<��Z$g�c�*7@���BD�@�N��C�՗�x��vM>�����Yc
 ���1��g�A�,Z����y�������Y{�Ԉ���������Y���Ȥ�����KJ��t (�2�v��Bh�Xg�pd�k�z��U݈Ϣ������~���lٺV��g�I� �֓�:"�sﴺ��QgQ���E^�)� �)���c�ch�h/������&k�;�4><�r�E�9���(�)��l"�-0��k�3������Z����r 5S��m�s��c'�x�H��C߶�Z����<�AW�J�����U����[��[����� ?��9�\,AXm4h�d�����w�1�e6K�u
�s(C�`�D�?���,���
�+�|�o5�Ah@sE�F���cZh_T>�Vf^ۚ�˳~g艔�{@5��E.@����9�1�I�R��^��8d��}��$�ϙ� �	���;;.�ؐŏFQ]��9n�zۜԮ��4.�`O��22|���+�F��um<�3��U��*�b�����������Z!j�{ݣ���[	&N9����; ��oҌ�;4�l�8�q�"[����q	�N������W���*��K#�F�Ol�Ge�Њ�}�p����"~+v/xy�+�7:;"�����Sz��%CH��63��(|�j��Q㤋4_>�[%��9�K/|�j�θ0�e�6��H���&_����s���ͧ��E4�+��=h�jru�K��Uy��'S5Ou��5�{X��E�qd��Ajt{]�@�_vn� .��׍�������=L��e��o��K<Q�+n)� '9�F��UFC UP�=,*D�o��� S&�]~��gA~��ۚ�s�l��!K{;&�T�r�
u�~/�`�Wt�i%~;1��`]ċ����R����j\�1���%l��J=����U$7(��^LfɅ���;}���pF*N�]�	��Q���M����.g�I��w
��xQ��-��kϾ��`K�^�IOqI�X�e���s#��"�/���I�^q�{��:r��8|`�j�)C��S+~��a@��$
U�T�Xu���C}�#��O|��hҫS-eZ���#��VqU�!$�ꁽ�Z�E����4+�J��) F��Rt�fԚ���S]yB���^ �m?��8&L1��lm���o����̖��#���1M��9��Y�Y$��C�����`u��E[P�9����t#7�D��25����N/��蘽�+"*���T�W�IC��f�8Y���JE�>�'����=(/fR٪b	n�ݧ[T��ʰ�5�$�&V�����#q-�ԓ�	�b��'i��MW��	5��7�ܫ�a7��8(�|qM!�����&R�����/�L�9���+�Xn���^H�4�QD'Z���T^O�r�g���ޭ<}l�5���q�_d�]�+�_�(��0w"�� �4J��]�=��e�s�̐�1Q�#$\���,8��8�����z��2x/f[G��#��޾�d5���9d��cp���8�$j2y����XA���]��Ek'��0۠#��S���>�h��T�d�h�eR�/E����uf�N`� Ǆ'������,x��Ȇ�dB"Xf�3C�pI~�e��~��q{�}ÿ�A��ׇ *y��9 g�59cS2R`���5)�;ꐑ�3���7Eo$`m�w|ړ�XR��&�^��8�<@�>i����,���g�92�����ba
6
fqX���־��I�*��
����g�T\n�N�V��2%�ˈ��"��h��&^�A�7J�rl�Nuʢ� ����Bc�Ev�G1�$���g�: T��V�D`C�br|fz�D'��9!�?|67���(���xKG|����v*��/겕�E�����e��*H���^x2G�������v�\��JU̠��C�?�mJ{R��� ��/4�`�����$��c7
K|2�4�@����Cxc�s��g���;)��e`A�����+cu�Y�,z&S⿿��	�kl'�o�\/���B6����b̏�~F(d¿���x-F)�f�D�F4ޙnvd��_��zg#1{�h�>�p�M��lV�S �|c���Ca�� CT�F�y�G��	���$���u�6���WI,��WWW�Ju�?rH< �{�F*dXFJ��� O�Y�(u ���q�;����*a�'ܻ;`/��t��,P8.���ysq�R�"ߥ5ߓK}�ͳ}~��"j���^
Ґ�^I�}�'�W����p.-)�(�Q^Y�<�BcƠ�@�e�rfzW1 t�Կ�PM���/�8.F��{V�q%)���T�8�F��"v�ѯx��1�,��M����	�:�!sɩ>y�RvoB�Ų:AH�������J���"�[}������~��#�$� ���iC�H�|S@P�E��zm�X$��U j�P'�ȏ8hi��TEx��$h�{-/����h��x��賩>�S7��Α����$�A'v�VL2���#�&L��tp����㵈���39~���������j彡�g.7N�7̠f�p��[���̮+�L�b�������J�uJ�Ӵ�{����D�����;��}�N�l��ػ+b|�#��F�Z�*��4���i��Z���q(�UlC� ?�dۅ�R�:�|�m!�s9/��Ʉ�g>�ÆIz��x�0��*lc�fie��&mAj3���O-I �h���U�h���1��+\�������+���6Fv���;�^z'�ϡ����V؋-�R/Q�v��H�q2z���5�wM�Y����yl(]#�������q�$(�oZVڃ��.�Τ�rc��
.�pd��h`#F�78��p�/ݠ9�L�e�Z�s,�oy�?P���׶o� jC	��6~d�&F���W��u{����`�Hq�mh�U����]�\R�c�ஶ�W���A����ٍ��ju�5i<���� �Z�Qb���ol�}���V�En�m�ka�O�'&I~9�3��nW��w��(<���紋À"�4q����x��qA��Ljݬ���Q�;��Z���mun�q���HJ���o΢_�>�!�,���v#���E;
�2j�X�ST�ѯO9�������'"�=�W�\G_#^�c��}�I�a�����ʔ�A���v� )�Nl����;���˙Krb{m�Z�^�o�J���BH�ʗS%&�P��4���I�u��5_c����Hvt��~�7LVX�9f��1��0�Pq�@�Bqd]�×_���W�����j��x�g��n��x�Tcx�ϕ��~�q(�y�'a�`ПT��O��j�!��qF�Y��	���۱q�`��Ķs�=����z�^�����mA�K�\�ymι�`��ɭ��j%����a�6��CE�CO<I�k_;n��{��8�fɴ\�bu�'���-��:����7Ҳs��b����=�0C|\�0���'x��9������'�����Kم��,ћ��]g���&���֘�`��<�&�5��M�OH54|�\�'0�� ����e�� =�p�t/�b5��WQ��N��������;��`���=�(�G>%�c߫j������>�ǡ�bƳ#��[��tK
�+lx�U7�����욖��T	"�-���\��TP:�1���X�Y�E�[/���in2��j,�v����'�8_Y_�G_�{����1�--��m�� /�xq��"�N�c���B���N���?���4y�� 8��5_���eW�֌3���A����ڋ�O�S�DJ���>�}5ʅ��\��|t޾�q�B�z��H���\���;m:�7��ec���/�R�$8���8����h���W#'��e��OK�zG���Gc{i�{�6��-��o�Q�����;��#;�T��0��өP��$RԪ�@�T8��ԝ(;Kվ�ʽ*Zܚ�֙G��iw�}D��]Dm��g��KŴ��0퐆���k��ʙkĈ_ӈ�_*I��(�+/G´���z�I��;v,�T�,��I#�D�=��EIĶmTjM���S
p�P�
��fil�dMM��6���?��x�r��W�3��洬�������	B�J�J;ނ{7鯳���;���:s�ߏ�P �8B_���r��������g�<}��F�>vRLƬ���k�|���ݶc�E��H��W+�N�0
�eλMw��4��+��������JQz�۲soe�����S�T������,�w��ia��̑����	9/,���1n�fh��~��y�%�xB�:%�Hg��:Z�<J�y�

pݾ��Ő��< �L%:��F�p��-��!w���j##�b;�e(5?�G>�U�7X_��cǩ4�"O:h���\M��Ǖ��O]���׳�]h'�q��L���y���ѣ�IA���{H_,s9CG�0Lr���A�\O�ɬ�s[.g��0�����uE��,��+H�^ݫ�/>*�{?4l�2m�Rx�W��
��9��^s9^+�U}7��QnLb �=se��Aٔ[�x�]W��J$�Z�g�����������A��ˠ�k��"� �hX��=�O���*�<���[�C��E�E q�b|��� f,���	f��W�j��8� �UȘ��U#��f�\��/�<���9(�FLO,����FE����,SMg]�e����k����s���S?�=l�k�`��VD�K�����ù9%y�� 65�N�V�Jݧ�zI��p�xoWgÐ��e�I��c�W=x�/�Bu5���b�rƒs�M��dr��rӅv$�e���l���i��P���f�C�s��k��n�	P[n��<ʎv�56eǒU(R�d��8�6�|�V�+���j�8�lnV�r��ܗ%�(ߐ�Կ�w2C{�b�>XlxVHYEB    ab24    1af0e���+!\�{�n\>�mWa�-v����d\�����Z�&�`s��
�����Ɓ�ɼ���gu�_���T> �a�Y;�/[�E��%���lr4��J���mCn����W�����O�̞��6U?�lT��(�}�8�x���@��r�m��	�C֖N2�L�Z<��S�r��:@�J+��I_�o I3�]87�����_p��W7������b$��_E����RK}p��)z������^p	L�1Y��-�mo͉zo���ͥ��r�����n0L��&3�iu2�= �cD��gP��	ZGlj�\��IC�V?���~X�h-_��$����KI=i���!pd`nl6؁�c@�oCj�� w|��?Ug��N���D��D9꤬/ԟ_лO �g�7��Y�m��"Q�ri+5D�^�!$>�� ��}��e����HW��ՁPP=齚�~�^���R��m˚��m�SI+��m�*���
��(�$Z�%����"oPX��ʷM\&�6?ðu�Ҫifq��wM%%Ʊ�p���ƊC޷c�@��#�P���w�J��9����-mk@�l��I�>Fb��Ѭ�;}��}���ۮ�f��;�|�¶8��O�i1i���ז -tA(�|u���T��~N��h�������Hg���R=�5���Al����9L��y��O�\4�M@�`'Ea�� �ia�vmF��x�7=]}9�ǚ��Ǟ}��-��XEy`2>f��/X)�.�g�h��O�3](D�N�t���s�g�LqΆ���t��W���U�)
o�pD����Bx*��k�Zv�ą1�X�����0~!��$�|z�F�U��&��r�8�)�?XLS��w���f�?�W��_r�2�A���;!;��e��*q���i3|I�Hq�#���fW���x%���4JI�I�s#��AR1��5��h��X�[�f��w ���ZymU-p.��]e� �S��~�ß�G�A<e�Ym�󫜰ͼo`�e)<��!Yx`�1.��Gdn~EZ�K]���"D ���S���gn�$Ny��5�\�(������\�_;�F�J��WK�"�"@�2�$a�m3�ҝ�,�Pn�a.�/��p@{f��,v��'���� ɶ��k��Y/=w��PnT6�Ś�:r������Q�(8�.�66i�X��W�![gysJ�)�)�տ��o���S��М�zne'eG��w�ΈU��	�U��ۥ,�zYvZ1�z��@hg��sL*KL���X����~���UL�r1�S�a��G��රǓd#nRF��(��ڿ�4ʓHf�H���3Y�U=����6;ޤt�zl/�k�O���'ޒ�5m2�S�ʹ{�^�Sb�.�a�խrC��UU����"M���q�Zhne�95$i�����W��O�\"�7��ES>��U��*��Y�ߺ��旎�3!�wUz�2�6�r�AG�\�H�W��3�0!�w�}�(. z�lq�q���,a��Gx"R/_F���D|��3�k `�lY���uB�f�Oq�����9~C��Lĩ��V��Um����=9�Z��ǈ_��6qq��h�BǍ)UT����F�jм [+��# g��O��taj��6��OCNZ6�`L}�0:����T߅W¼��y7��e�S �g)��7ŋ��q�;�|�����+�|��$�CAw�7̄M=���}��I�6��w�FL̗�L~Q��Hg&Z�)��f�D�R�98i�T���܋��F�j}�/���YN��V����k	�a�K��V�B�d�J��\�Y!fgQ��Ё��쩗f�l�0�s�7��5���U�V�Gd��_��������2���"h���А+�u��wAt��{� ~-o&�����x]7��:��K*�$��|F��
縮�p��.���\��@�& ���i)Gw�� v�a=�m�+8��+����Iv� �ؼ��.%��h�(T�ţYu��e����,Ɛ�:T+�>��m�r�:&v�>�?�K���F�w[	[�����YV��{��~P#_�8c�����X�x�X���@���O��el��tz��:B�,B_s�HI�Q�o����&�ꃕ<���K���]`����@q)O0��&�u�6��>������k��Jz���r�W	e�@�]Z�,��HX<��W�f1�8�����#�r�$� +��X;Dt�3���_�*vt���|5iH�OQ#��]��c\6οl��tϑ��h�iS��D}�,�����]F��|�f��ˡa�h�u�2�Q�����a	#h�h(�'�nu=��	*E���r�3xgC�1C���t�)!yȱ*H}�c�Ky�M�goJ�l���5�������ӊR�ڣ��ר��M���g�@�d��8�6*4LG�|^6[��u�,��W��d�Y����t8��I}�P�N�S2&H�Ʌ��L��]�);JF���x�E`ԁd���qr��,�K��a���CE����pC�'RY�"�[���<�� �����-S9�ӟ�N��*�T��K��;v�aeF2"0cU�?��C��&Ob��2F�:*�������5äe`ߜ�~`d��ƍ���w�[�U���E���_���A�m���MĿ�W�a��HUo��>dę&�,��m9U�^z�1x�p�Wd$
�D�qΌ��ݫ����@�
�,�P�sd�x������k����+\7��W9��g���㠈��e�E���.����B�S��gNa�V�z�`�a�{3(������<���uF�zcI���Z"��-��*�*B��u��r���r���&�}�v%S6(.O�A����s�-v�q+P͈�)P�xPa b�z�$5�1�-���-E*dt鿤>),��+`����.w6�����d�nZ��~|xΐ/�����Ğ��kl�C-����n�Cą��	�����F�k�Q���_{]�H�o�G���������U�XJ�����4�+V��m�;�kF����"F���؍x�(6� W_��Zw��s����א5�MYLD�)��|�^4�A��!�b�*��۵�Ek
��}��Uir�H)^�w�1/�Sø�@／��6���.���<��0$�Nl%�yh���L��M<Ć!�2��r���
�ʊ��J�r=ǘ��}b�H�R�ד�s�fHW��"D�nX��E��k�	W�U�i����iՈOz���Y������Z����f��J�=5a�
OO��\~
!�Z�^�g�8=�^�-�����D�G�M�]1��a��8L"�u�yut�J�c�1��s&-���8Jy��p�
��	�p
yấ�@zb�ݑ��\��C�����[�b�|e�'��9��0��AK��n�nqz�~U�,b`��C�ݫ<�~�㖅�vE�^`�xR���2x���@����9���B����ܞ�ꨍ�+����+�&�v�_׶f��l��9�j���-e*]..�?u��ŷ+m���[���D�_).Jp}�Ѿw/��;��"�E��Uwv����z��Q���渗�Q��:��H]�'?��h�ru:�kA���R�d]�Q~���-q׭��r�f��e/z�{]��6�4�7��-�?b ���l��쓽y^sb���WN8���:���
ǙAh@j�\�2>��~��2�O����V��<�co�O	vt֙+�命���I<#�_����rY�Ϻ��Z丹�*y�ؿt=?�o�߮'�wѮ0�:x:��ÝL|hH��i�P�Wb�n	�J�����[�9�:�p�B4�=�'�#�'#	"v����"���Bl�yx������"�8
���MQQ��1]X��d�u�Pg�.$H�F�̧ �^8H��u7ǟ ց�hkQVI��4$yV���/�.��������Z{,���<w��Ԧ��������n�:�"tA��|	��j�M�Td��>Ø�.9���6R,���Co�C�)a-��Q%�Hk��8Vb/���l4�:ގ�j��2#{@����H�lF�h<s�|l9޲�I�>F�2�}Wg�-��p��Q��8׏�n*��'� Q��h%����r�]~Z����To���WjUa%~�[���M�PP�E��ɣ�����k�]�o��	9L3���5�i��S[����-���!CpҸײ���ϸ.i1x�{�롲�Q$��q�<�د8�{;�KF3e�f	�	�~	)1�W6d^���8W�/&{��ǕD��y�G�TnU��ӫu+3��#�LY�pd��� У��&]o���p|�h��8����H��[Q/E;~��`�R*�w�:H�Af\3�%�e�E� �����6�!����eꕥ[�}�O(�O��Y�$'�&�S�{����4ˈ��J�d�5�Gv�+ S_��������gkG��@<�QW�^c�ȮE,�H�����Iي��$��ۖ����PME����X��Q8��ћ�eeI�@��֤H[�O��R�=�O ����X/QP�NE��W�^��Ω�(Fi �a�|'G)�ei˹��D
w�U��߶����*==���v$�WX\w����"��T�і��#����5Jg#-��m3��\L����gI�1þ~�X��S"�(����.�&����Z� Bz�jަ�����	 qJ�:�G��'U����/���a:_S��!ӦZŔy���<��?�җE��w�@ጡ������J���3Xu��E*�}޹��3T�L��5�J���~���n�_$_�u�yje;�R�z�o�Ģ��V./<ɂ��P����43���W��Zuʭ�������a�^b�;�[7` 	�I�g� "}�d�$�L����������y>�r�z��s��3<ֆ�`��'�#V�5~\]�h�WE�th�K h�8��T�V(Ëk��mW�^"M�#N����l?�����/ˑ[	�ݤ�����Ő2|�I8p���##�a�naU�i��ؠr�����.v���]�� ^&y-���^-}p��#֏kU�`�������և�/rX̃���HSީ��P��.�INJ۾��������Ѹ��Q@�!��5�<��6��K�9�8������O�#ҵ�	6�F`�9��㾫�e�I�E�d����ɺ��R�9��y��L@�42��7��Ug�q��.��z_���Q�7+��w(����L����Q
�z�.*z�U�,��&��h��5���`)�pF͜,� �׹��~Q�x��� r�W�QP�&j_eI��f� ��D6tf�0�U�/��w����� J��9Ck�9S�"����	��X���W�4�6Nc.�v�)ø�ZDRM�)1��ee�U�d�*n��m��ϵ>���p�R��:RF2��U]�UMv10� =2g��]E�>�U�.����� ���,��Ls%b�� D���,Aլ�/�D3r���N1 �)�v�v���/��C%�����@3���8�(�j�=kW��L"�'���JA`��,>�!�$��~Rp&��� U�	N�@8!O����ɒ�p��}� H(��/ܐ1�@t4E��C/"H#����}Z���X
�قq���7�S�?�P����kO6U\�ݱ��v�s�cz*@͘��6�&gN�u>���ޜA��l�C׊f8��tSr���~��;P�V�|��c�����:a:��=c �Sq"Ϲq �'3F�T`F2���I�ֻ�t��rz�F���\;���J9����O�"��0��̹$�,�`�d)C ���������sa68�]6�Ow*�BB��&pQ�I蚬��X����rq`=#� ?H�q��2��U8����X��bG����:�S@/��;��/��m���ҋ�7���0��̷8yV1�9��^G:��*�,k4D��@[�:�x�����, V����:w��\v�VR6���	t�.k���Y���n:=�'t_�0J7-����V���5��rكn���bf1 O���f�Xiv���<�7� ���O�Y[����?�$���٫Q"H�בl\�� /�$���G� ��)�\v��u�4 �ޜqC~�����Ѫ��B	,q�~�|=!�dm#�:WD�����pTϝ}�.�)0�������88�N��ėZ��A�'���P����h9-Qָ|��ֻ�Ȼ{��YS�.=��v:�h"V v)�᣽�i���\�}%ᇽ���P�V/�a�)������$�ӕ;g����F�O��Ju���1��R;њ�Ȼ�b�^�'l���Bޙ�.��b�t�f��֋��Dx�??:����`�]4��\T�A��y&���^���Q��'6b��,��n���Lz*w�������O��@�U�s�����nR�{���m�<�A�r 1�ӟ>{����<0�@րH(�C.:-�m�$�DW#@����dJԌ,�f�~�7���Q�����,IܹkFHG.�#�ء��i(�qF��PQ�8�������0�F^઺Ǡux�U�O���۬ӡ�H�#��8ע����o&���%��ծ����X���T:3O���D#�� \���DXL4���'��y�w�TY,_�?�`�~�[� ���6fZҔ��c�&�8��"�s.5�Xs��Vp�~�Ø�,�m�yP��u
�[D`�ɥ���8�}u�1RCU��q�1:8�6�]��V�����-ڄNg���۲�