XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���6��T�\Oٷ:�w��%�3��<�C^�����]����I�?���GJip�3LdF�{6�kcr�sz��r��Ü��|o0�}�"���i�H�@Z˖�L�
���2��?G�<��fJTɨ����M����8hR۶��ffT�����\δ���
_I�u� p#uoZs�����m���H���u�^���k��:��/�ZR���q 9¿K	0�Q��6�����Jpe�U���=S��	�
�{�Ijlo2^4V�(�7_��-&M(�5��8��9@������#kvZ�������2Ǯ�����d0���v,w���/E�?�����$�� (L�i�d�|J
�_.�O	�$�_�����E47�wx�<��ly��H���f��aIJ��.�{���Z\�
�G���9���lu|��G���m��C�-	�&F���<�嶒F[�EŎ�S������ʙ�n��{ա��A$SjЄ{3�	�"�[��@$�Q*�`�h�xD�;`k��2�~M0�Sx�<�Q������d�ŋ����a����Gp����G�Dwx5zo
�� ���g35WUo�皤�c�gP�Yh�K�s�1��L����|��X{w�b]g�C2"���n6n��y�%�lW� ��N~�a{�
�4Z����� ��iW[��:�v��s�1W',�ͮzct�T��,Z��8Y��s&sa$�a���D:c����nG5x�E^Ԅ~��%�j��y���l�6u��hXlxVHYEB    22a1     9b0Y�F"��*������rA�h)����mz��GG����$ ^��3m$�w�~��/����S��UH�uW���&���v��@�g�
���WQ)ǡ&�k��x1�3bʟ��װ�Ͱ����[|U2���Z�ۜ��,cԐ}�'^�a"^���E�B�E��rFm癛�A���5K�bF}[�qK9�ϔz�_@����,�#�B��[�:��K&�F;W���"�x�vh�َ����c�]ك�����;�/��Q�@?G5��o�?��D���|b�.����	��"[�S��<�DŽz�]�Px��0�"Z[�um{�Kee�W*��-=+��wy��a]VO\U�^0Q0ܛ��b;|:�/Q9��-���X�q@�v�Qi	]�\Q�A��x�)J΀^e}�
9D��&!�k'{Ё����U/��PZg��l�@��m)�6P'�u$0�<ik�^�􁫋���+]����
��1�@����t
��0Uf��A"e�����r�� ���'�=+@���}��|iɺ]ҋ��S�GRt��r'�ް~���*d5��@�Gz�le�S1���Ǥ �DD�d�̫�+fP�'.�"z�F	��>N�FK����ʪ�����M<a���Pb��Q����5ݥ�kK���]�U��$�(��ڥ��٭�2�:�f�w2Mc#P K���/��y��h���%G������?~B%�rX��U�^�$.��M6dg�2"��<|�.s���=1�qb,oROW�sf�SaCZ'�U��A"§խB%v���T�zJ��ju��h�C�#�d�Fw��
$S_���$��#7ѿ[�r��4��pȧ5��f������V����+��S%'kI�'rH.�z��1q�H�~��(_YGG��6]GV8������>�WQ�&�������J�k#�l���TI�,co8�7wwJ��|	��V��A���e7V��ҊO�Y�W��V�kD(��DM
ڧN��y7aF�P@� 9.֫��a�53.{�#HYɜ� e��X�.��IjxZ�V!�P^dO��*`�I.ښ�ۢ�;��>a=\�,1I	�y~���� �T��l�)e�O���O�@-�)3ӿH&�E׍V��p�Y�(��E������ц�x���Kѧ�y�
X�xH�Oښ�� G����	3��8���
E
/��Ţ̰z<��[t��D��?R<��DVyt���T~^�ܝ>�w�rr�|h�箎�C,_[��p��O��[V���Cz}�i��uU[�RFz��%��ee_�����2t�J�AQ�q(�54����<V}w��q�$��p �@�w������*e�:U�8h"J�(�ǔ�*7�1�Q��݇u���HK��z�4k"���?�}?� ��[1	fV><
©���v�`)�o�H�P��,��#�CQ�&ӆ���#r1�t��*}�;����\X͋��W>H2*H4Ik�4}N
����U��ђ�Q�k|Eߴ�2E��w���bsȻ���P]��Kp�Rs'�5�πDaT���{#b\�R�Kj�0�~Vhߐ�����Rl�ڲ�&w�)�Fv�'X*^u{�~��zr�MOu��c0�i�R��%�Djz.�tB�H�2|�;r���L�=U�
&!�y�}t�u��e^̽}l�hE�K!��X6�n7�"1��9�FJ��q,��ΐm��4�/� !������Q��[)��V]��f�dQC9/���#��p�db�۸],n�ҋ^H!O�+p��vVG�2C�B9�WcW����Ր��	�����#C�-n,���(���ؘ�猩
а��ޡ�Q���'����U�k,?ɀ5d�#͡3:�O�=�H����A4���8=�m�و�ӷRw����mF��3�ݷ��u(��e��UU52����I�ϡ)��4�4��!�м��!�y�&+��w�5�������.?��'`�I)�+�m�	�]�������X�z��JK�T�Z��7]2ك���d�����6�zy�.
g@�܏,��׫lD�Z���]o+�O�xSA�RR��T>��6��]�NK�~L�E�6�V�V������:?x���>��E-k��c� �3-X����\"�-j7�1���e!��4�����h�ݟ�oP;?�F|c��p����o\ך|�Bqݧ�'F�eL��/�%��7ީÏd�DUr��'-io��O{C����ur1cqlw�Aaa����0�)q���sH̑g�{�\D���>� ���*��m�_ٚX���f]�]�f�X8���]#7x���.���S��fHC�{%&��d�erD���x{IUd�����pcZr��1�[����
���n��}�ʈ��M�����k6p�A�7]��U���"��̈́y�L˰�B�V�B�b���%
����^�"��m-EZt�����w�/���a�gf`Hhi��F.����w�n(�DKa_�