XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�v�r	�9�闑z@)����vQ<{]�֗���V.؛~(���/k
[p�k���;�����님���8�
��t�v�wL�)n���%A�=%D0D��
Ò1��ۚ9,�g\�c���Xܛ������j?f�MR蔄i �<��a-�Jn�y��:��-,Sͦ�y��s�Fͻ:;ʅɮd��nʢ=�p�^�`L�)�"d���=�ia@�-��P>6V�5���D��Fx�n�LoRq�,txC ���4jkpz<�	�]|Y���l$��Z��i�,r��	0�oh�y�䎸��Ӆ�d��P͢K'�	K	��=�5*XAa/5��'�+sNc;�>U(6;<�=�M�ha��g�F<}]����at��k!����w9&��*ʖ��ۤ#^rY��{A>�,�1u�\K/�[�K�%��#;ncJ}�'ދ&{�1-	�����/EaEUӦ�3�Mͼo�w�dԑf>�V��3Jn=d���^�0�����jCO�Bʻ��s:\���y�ѡ���n���]�ԸSu&F����z8D�x��������j��u�aoOn�@��Þ
L~�
����Mx��<Z�ހ_�-��(GQZ���=��0�1;��$�94��ǎ��[��@B�tS,��E��ŅE�`�/TA���K	���uu��v���0��yA���5L����0�M��tl�s��Y����ƏA�<`�g�*�Kغ5�<G��b>�r�O&��r��lbbXlxVHYEB    1e87     a50 .\���\�w�G�ip��O}aS�����b��tm���r7�[���eX�KOX�ʩ�ne�)* ���A"���ڗ	��<���w��+�S�ʥ�	_�<�&m�)7��=kv
V%�Jd�"!�G4���۝I��MՅNG����"xzn��o'C]��A����6�����s�#N�).���,�`r��/�ϟ��F9�Ws�
���WU�r�����H�;�i���~���Єqafl��YQ�O
KIp`�A�'�uI�@o�$����-�1��.86����J��J�5E֣l��n�� ���D��Em����8���=�C��/!"vgL��62Ʋ@�1	�ޜ�˴u���F�]v�U��k��Nx�P4=O�����~�`���������B�u�yb��v5O%�����%��:$���	��"��D�v*�����Oq�%�㎽�dh�I��\:�M�ٲ��'���d�mɏW٧Mp����恗���Mֹ�ҧM�9��:�6IpY�t�|  �3��%�f�G���,��``>;���\�K����4l���Z�~Rǘ�ʖ�
�m}����Y}�(�3.�,l�w`��gw�n�|�����@���rs=3qO[��_e�Zd_WMu����X��o���L�AsxR}!��V�{� ��>�Z�ܖ�<���N�O��tdf�I����Z��[ŏn`''���>z<+QkdM�&��vt���xY�t	�{.�D9:+���!����\N�^
.�3�����!����RL@(�h|@%�q�3������|�В"��6���_�
��`lW�6���.��CT"+'�mTQ߹���::N�x:�Ϊ��p�ǀ��-�b�em���C1�*,_�,�M�ݼ!8bR{���d��W�ʜ@:p���(L������=w����� U�bm'ז����@��2�:�U}�θ�/j�c�5�r�%�'�`�h���Nsxi��pʤ(Y�(�!����A����:��-�,|��1�+�pks�Z�*�ͨϷ��0#��Z�O�u~j�ǧ�C�=Kj��<u�)Wv`���ߖ�PjcW��[la�0�B��� :ȩ��j}��d�\K%:�g$2x��iL��r�j��:'X �N�r)5��1)�*�f�0n&@�w���u��y�KǢ�}�r��C
�a5�8���F$#�����������+h�e�3�4�L����
������ۺL��i��������Ɠ!���?��(w�#�s7�˫)���h%ޢ-�M3|f=�ƒ��S��N�רԠ4�Tu�8ϙ�V�/���v�KAlxw��j$/eЋY匪����%1�,��7�u��L�YH'W&���j;ї�K���dw]3�u��E��h8Gt��N�.T��^U��(��k�yC����iI�8v���h-���=j���B�믛*�#<ڪy&L1erp��=�'WKŞ{5��~Y+�o�81-1
JȽO���HP�ꃷK?zD#�U���#b$�`U����O��*�oT��R5?ja���jk����T�g"E"���v/�3Բ*�bV_��1����O���aܧ+7Ju���'6[�	���C�N�ނ�I�H:V#D�: 9aYQ���]�5I�� $So�����P�l�!Gs,?�!���-�-��ȼ�az��2F�𦩴?�%�W%]�D����Ͻ��j�-�����ǃ�5���s�͘�e�졯ĺ��Z�=zt8ēؕ�U��3�bh<���,Lp�k@ۃ>��&+�9�H�4�{I���@	ti��5����SS��.>������Gb�,Ř����9l<���|=/~
�:��CG�������hz�ʒ�פ.�d�M<�l*��цE�4G_V9y3}�<�i 5?�+_-�g�*���_�Sv�g��1;�y9c3���|C�A(H��q%��a<�	�����m�	ȸ��mc�m���(�p��?���]�y!����� ,k��Ӣc1A���3�ջN����� �o�����b��=�/�џ���^8�@m���Y�~ϑD�R�5���b  =ޏ�Ɉ�mPT#j��e��]��Wq��O����@V&Jji
�뺭�(�l�N�!g��d����3D`Kf�ɶ��a�B��m㌩2�S�V�����E�A?�ե&��a���f��mB<������4N6���q�Z+C�x���	���W������<N�W�/�Ğa�
��-����M��56�G�d�����m�n��uҡ%c"�ۢw�1j�j;H-��3E7��$�(@����2_�K]�]�4��3�,�\�b��Xk&��r섯q/����hQR�%��.�&�;�k҇�!���HG,�dkQಯ�����e[�����j$]���9=?�@�i3�K"8B7�MVf��Y�����T������6ί
9�ɿ��m�u���q�Ɨ�Zt��s�2����X
� ��%���/���@�YU�O�'�)ώ��r��_���Uq���� �x�Zm��I꼡�+[u
{���?�ƽ�mq% �h�#7��7^�I�����Đ�TO�#�� Ƙ���^To[�2
v��M�9���K 