XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?�xr)=��yv<�q�@< >I�}YF��$���p�#���X�7_��/��4�2ߴ=���\h���3��|�+sN�.E#�,�2��1�b��,Bh��B�{w+�E�)މ��k��7Z�-漃|22d��k�����4���A�[�9���L҄�8��y��\[p>��3؉��Ͷo>���>A�J��!�!�k?fPf��9�&j.�)C��ԁDY��:Ǧ��R�	�qX�T����6M�F>��j�� �|�uP��{���Uݏ+�v3W��<˶
������e-���PҚ�{9JD��DȺ�m��T2�K.��.��ΨZ!gU {���뢔�U�bX�yq�V*��r���m���]f;�U^p���I ����gg\P�L��nc~$���A�̧TiZ{�J͓��@+������?�3���8�����rT�̶�/��Pڷ졒�5O 6�Ҙ�D�/'�U�r�t���JOb�m���)�n������$+�w�X�%�~z�l|��ɗ"6ڑy����S�7m+uw���v�R�c����--����1/��'���� ;4W��ŷ��G<�.w��\7&6�L ���3�c^��u��a�/���coT7�%,*	 �(�����7 :�#{��{���b��dG�!�`���v�wM�4/�h�џ��F��X� �xb��d�MqY"��8�^���q�9M�o�-M;YM��N榒����'�����<1�l�XlxVHYEB    1b40     940s��vй��c\Xh�W�-o��@G'/��g"!����6�M0����d������jϧcx��V}y{纡��8��A�O�'�ZN+�t��V��>p6e���ZVud�ӹ���#�p�-�p��˝��3~��S }8����Q�酔IE�4iZ�Q�'���*T�_Y`b�Ub����?FK���N�Z��0L INf��f�f3�,��.Ne��zY$���/]����G�<�hw��z���`�a�yuF���=�A�cq5@���B�*�8�
`h�}���z�����C�2C���c���
�I��R,��tn�x�^�y9j�c>��"pF΢0c�8���B��"�+��K�ǚ���v	ٻr�_"���y"A�V�O��-��]��nk����lJ;�袆�����:ꃆ[t<���*�:���|u"/�ۉ��~����?9C7�ڤ81�(M�R����6�_����p��׿��Bt$�*
����0��f��iW���&�o�Lִ�\�'TT�1��)f�B�dO>�b�g:%�9�M�ʓ�����%�5ݑ��I��U���=<yHG��tV�P~����`�Z.8;�K�!���wJ�������_m-�l�C����M/^�[O�y��4j��u�O���`M�l�y"n8��~g��n����%���p?�����0[��}#r�b �CW�	#/~�O]F��:��U{y��Yl�q���M�e��d|�<y��tЉ�:[<������ѱ.� ��x&�i���mPv�g�؟x�A!9��t��d���Q&�H���b8L�4��VG���1{���[���\�&��-��p�7u]��Ӏ�IP��M�μ�7��g�M��ų���R,�J�F�KC������
ec���tDJ����/.r�b�^,aO�PH���G��ks��R�M��ꇈ/o��zrJ��%�K��P��1�U�}���ܢ`8Ё�ʦ��$���v�zIoj��h�	1[3�t�y?'�O�Dh�g@��s"����#��Nl�VN%� >5��#Q	HݩCs@��s�����hw۪E1�p�oC:�r�B�؈y����P������\�A��N��B��v����:XE���㠸��[;8(ׯ��v���bS4�6�W~C�.I΁d;J��mXR�CW��!R�X�y�v�Ygfտ��OI��p�'�"I����_�����#X��g#�5P(�X���|�=j</Zlw}��ܾ��L)*ܖ5��2��AIXT�S�qХ���(^bp��f�#��T�8�RZ��0F��K2�RzK�'�?�lu��ݖ�G�a�E6j�T��i��ի�(%q��M�m1�$E��l�9Y�=����c�����K�;�xZ$��H�#��4���</���r����:�a�$]ؑ�O��1ݯ�j�n�O���G���o�?g����N��o᷈E��U��Ԡ!֖O���⪱P���zj]yI^KJe�s��Q����|���Y'��H7�u�h��e��u�xe�D�?Cbv�ā}�{�'���W]�"}&U�'�����f=?ɔ0(񗋀z����X-(�����xv��8�,���j�z��@?��!�Ƌ�U8A1�>_���t����sAEGzT.����LO��b���if��=h��E�O���eZ�����&�����×t�����\I�4��Y5���ݾ���^�)�$(�+�Ų����7�{EU����h=���]�<?ė���sD��W����w�]�ۡM���q�\C��F��M��m��w�W֧��r� ��5S�"4��69�m$�36]��h��c1�Z�!�I=*�N��J��/����GF��*ï�Ү�+�8Pתi4hQFG������4qܤ>,S�w ?�{i��D��"Bq��ׄ]ד��<�Q0�/_�����] �������x|�f� h�������` :j7	��WQ�䚃h�ʤI/z�7�!����rI$�V3�2L�d���B�4(�2t��� ��Y{
w�}��2����2�{�����D�<	�T�fLP�w}/K�Fz�k?�t�$��g"LaVjA��|��[{p�}!wӵ�\wW+(�JCsd���b�Fhx���\>�~��7�vbq&��c!�O�UZ�l^c>���R>�^0Y��qZ�5�i���3q��*�t��h7��oI��	����<[��5�J��L��z���ϱ0@��dNb`�k/R�]}kp��e�����&�H�
�S�nv��{�rIr��Վ��1�Pڷ�l{/9�U�&$4��J!ObU�R���S�V:<�g�