XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��GGt5�S4��9�����գ��芖��:�@��;T���V2�jӈE��&�7��9�E;G�:߭���=�a ?@龎���D�0x����0hJ�}�nJR=�w��N���EJ~�i���@�7�?�ݠ��BH��	*5$�v𘱑W4���h��G�H`-�6SK��h��v����'�@��"7��=�w|d#-��&����Ӱ��#Ӕ.K�1_�3	��a��T|�v���L��ˮ���������n���~�#Mμ
������/K�O�oo��8��!	�����t��?���
�]�;�w�@z�_.��)wxc]b^ĩ��_(�;��0{�J���PȋS-{��$�b���5�lSc�����Ӡ�r~�΀Aq���e���`���=}j+ܾ`��I�')�ڧ����*Тsl��g~jd�B�qp�"��(݃:���Zז�cA1ĵ'R�t�Ǜ�����L�Ң ����&-�=\�yF��K3�#���R�#|H*���4��@��$$�O�x:�Ž���M���g�g ͝3��|م�D�ا�h��N�f(\ӕ=����kǧ1[�;F������_��v�3��
��b�b0���"5Ჵ�F�Ӷ�-��u����m��ER�}'H�.��I �V�Л�����`�3�"1a��@8e�55B=�������j}��5�2�jY֝j�$�;�U0R_MK�� Qș��퇋�������"�8���iXlxVHYEB    2a18     bd0k�5��-NG���Fï��E�� ���o�{��y��߄���2���9T�'=d���h.1$�I2����@���G�/̒�T��f��0�ꝅk�^x���P�#�n�4,����,�8<{^ٔ@U�-���a���#'�;T�CT~ڞ��,�v������o��G�x.�.j.��(V�8��Uj+%�r�1��	�\N�s�,�����:� ����,0�N[x���|J�_�PX����y҂�H�����i��gy��TYq�p���!���͉�z6�ol�m^=��Z@�W�ص������:�k�{�!s/�̜�H�в~�L �B�(^���|��\��wfP;�&��������g1�>
D��t�&-��~<_�ǰ�	�n��R��m� DPi_��t���FIf�&%��͓�bعI�$@c측��������i]/�r�L�6lk��wc�����򏀥�X9K�(6���'��6l��Sa�&Y@G�Z��B�-z����\���Ȗ���/U�;H,�A͉�@e@Nx K�"�=�e��vpŐ����=U�H^Y��bGíp2�:G�z�G���H��=Ol�W���c��'$픓�;�ivm?v������=�E�ҵw�ԯ	Ao�}Ǫ1�akT!�M�_���������`+/	�^�yM�9(]n,������ئW�si�x��\y�1�4ޯs�Frq5B �,bX_7���Y��F̝֊�l��J$��|����f�)*E���`�˪��OT������^Q����+�۷a"z�LԻ�o��W�0(F[A��w�n|I5B5�]/<m�м;
�Y4�������O�_���l�?�o�y�3��=<��b>�wb���e��HmX��܈â`z
�E����h�#\�G�� #�xL�p��Z��5���׸%o���%�%�����ϴ����e�+ ��{��G�����8P%o�\<�k

��6���{�B%w�{���~��rḴD�gޜ���VI�2�J���<RI˄��M� 0����IxfTF��%����Ha�"U����SXh��@��-n��]�:>c����iLF����a���r���!iBz���q�N�O��-������b7���|ڐz�ڱ��g2���!����E,�U��"
.��Q��/L���C
+*��t��׎jp������f��� �m��ja�C���������.e���>�3�I�Ƙ�-I�xKF���Q��{7��тL=��m,Mm�E "���k���h�ϭ�B�$)I��.l�m�(��Cf�N%���ԯs厹t(;��?�K*��-�F=��i�(P4^�,�����JN��˗��!G��+TG��U��Y��L�Ue��R�U�:i�y?`]5�$��!�#F�*E�]�M6	���l2T��lEZ��s�ÇH=
1)���~l6ʺ�<L ,L<0F1�y���G}t��J�	K��{i�c��a�A<�؝�zEf)4���9w��ca.����c3r���09��0������<�Xn8��,A`_�Cy�+��:B���_vYx	9d&֛�AAH?����*����<����y�L�$�_��Y��x����N��W�B	?���<׹|����$$=��.�ؤ���iq.��ow���
]8A�
� �P`��;Rܫ�% ~�s'V٦�-#%��"��s���Bz�N<��xr�8������}���V�pEU��_����֤��BFNL"7�݆c�����[J��F?� �}�|���aٵb�|;u%t�գ�^���,��(藿?�b����N�@|dK�	 e����$ܱÊ�᤟��fHޭ�y��K������U��Z�>�Aޚ�ts��^#��_1�Hq��*���� �S<� b�O��v��X�VE,��{�d��e�ݟ�e
>!o�h�}&�wK�.y��%�<�KJZr'�z!��Je�.�Y�wKw
�h�����q���`�	�H�eu���c�d@
a�	����)G7�e���� �G���F"����b�K����W��a�XK��z��yG���{�-^��+��WD�nD� SQH����<W��S���-�s��Z|��� �[fL��nT����w�Q�T1�]?�'/�wYfo�>R�@Q S� ]���2Ѽq�� �ڝ�p|�-"�ޏ�Q$kw��ei���r�B*_��2��ߑzw�Х�9��Cԏ���pM��C������G�Ƽ��(|ꢈ�7�bOF"%<Q�E��V����!�Cb�H���8O:���/�/������ꄐ�L��Ԭ�jF��#�����y�*x��`ʞ]�T�̊�f�d�s�J�V���C뚔����g��/������f=y<��9�XJK�圶pE�N���}�����$�v�j�j%�R�.�w��@��XO8�]�:U����)z��Y!��uE�����;�Ǟ2)��v���z���J8����g�<�Z#w��J��Cp;1F�H���������N9�Q�e�P�qo���j^4;�hH������8;�����K���w���.;IL�p)أ��[�^�w�|(_��pC�G��8EC��-,X�*eNd��$��S�Tx3� �xv�B�a�6_e7���%P�#�\D)��ޣ-6D��(���������%Ez�4�����)*V�z��NL�r柮�|͡�_�8r��Ǔ$�XP�IyWSm��>fij�-�裤��N@��Y�e��<y�[؉#n�R����"X�ܮ�A���i�� ���P��-3��
G��݊�W,O:j�Z1�(Y��g���nU��Q��2��s�1�b~sn���hB�(Jv�W��9�R��"��Fza8���23ج�-[B%�Nc��6��I�����|���_��s���Nk�3KF�NT�M�(��s3�(�a�3W�Ks�����/�Z�s�NL!W�k