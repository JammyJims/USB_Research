XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kP8� "d��x�*o�6_p�������U�Wyߤ^Cu㵱�w�o�!U���a����ȑ��0�����6Dӎ:݊���Th��|i=�uL�8y�<����U��
8�P㳎MBap�Si�#Ok�\1d]
�}�����R�F�P����_0ٖ0�Y��2�r����~_�s��x�c��((�̅m��% ��S-:�{Y��8��pϷ �;O�=�3%ٛ)x�]��{��ɐ��П�}B�f2��2��^�M
D!�#�WQ��p���=�;��`(�ST
O��G�_�c�|�v��f�/.�S��L@�K�	4zX���'m���l ��|�Eod��N�঑/5�����kQ�jM�Zo`�!iʀ	�O����*Y�!�?�Xn�/`<q�]� �4�P�ܳ��~�����=���K%�	�+Y(7�}��)j�^Uu����WN%�	R���¦����[�C/��KGb�F��!Y�=�mcЇ���Y#�ľ�3��>����v�˛l�R7��c�$eMO�=3m]E����gÛ�@(�i6�T��/dLa��s`O*�iP�C�G{0\�����K]�h��@|#Dq5�*�^�d�#��jN/D���jx���ӌ�I��R��	Y��s��Mt�t@�����*�r������ix�?l=�x��,�|l�V,��5��h]cD�I�����b���lP�lV�j�PJ�B�\P8��iX�=�Y��b-��e`m����=��ɏX�� 6XlxVHYEB    5378    10b0G�����`V4M�#��d$wx.20G��";P�_��8p�Ť���a�#�����#c��e}���χ�t�__�4�o]���`�W/
�B�N`��+Q��4i�L�~���u||k*����*@o���H�g�i�<ۥM$<a0z����ʓ\#/KQCCش�<������/c؊��`ޱ�u��)Jo��a�
þS) �do ��b���	j'�7�U�c�6�(���Ңο����j�]`���!\�9v�zR�7��Ra#�Q�|�Y�	am:�H���q�4��Ϥ.��������V���_�2 �O뮿���|�0�޶tc("(��0�� �$ʬ|��Dѱs���ә'�Ƶg�;�����_��w<@&�j+�5*i��+ Hwq���Nla��y^���!�j�Ts��=��g�Id�<�"�=@�]�T��T'm�IZ���T����ۅt�N��硂�S�_�g�ֺ �q3��3�~�Α\�qC	c���)���4�e�ܱ�&�4"�N�������w�+i�|���/o��-��Z�4L���D@�7���lX��&�FGO�$�B�h7"����u�o���b�E�MN��3�υ@m�����S�ˮSٖ�誢R����Ño�n�cV ����6�֬11�u
uP8����kn��H�c�-��gc�g�>��'��cx�]�ڪf���K
KͰI���֒5�s>:�������wZ��7�5?�cU�+�c��u�o'�И3e-x��LXv~����ɰ"�3:��>��
�ü3�l��_E�X�|G�"�X˒��J��6��Z��^���,[��e"�ͅvD�{.�����6�1L�ph�}qf ,�=���PVWR���;��]B�Ґ��ű��SEt-����ǐb5�
	Y⚁����R�]О����	�U���8�bY[;�R_3�D�s~�r�k�����w�#;���8��|�n�^:p��?�/[E�In�|XE������BӠ���W��_�Z9H�<�A���}٢m{Lz���E�	�%��ɼ�9�)��阚_Pb�]�|Kה�d�6��7���e�~)����u}+]��/0ٔ�WK�O�S2X?��,=C����Y$�Lm7G�����C���?zn�%��"�0�:w��-Ak0k�8?'c�����T�iHW��*NE߱�}�$,́��#!ܳ�v��/� T��s)��B���"�Xb?Q
����������)&����NJ�.2ObT�6]��&��	X�/��s㉕ <�!��Zຉ���,���n�p>��[h>Rj������e��2���݃#"+����V_?�W�A��E�o_\��|�<��xϰ$�-:jR����$"1��6M��Za�7z̠.�zޏ�Y1lI`%��E9d��$�ö�G#�hmq�]���Y���b[�!�Lp�����z�%�6���l&��q,�7U�"����z��po�ܻ͝��w�Ȫ��IL��a]�>��ђfs��(C���o$d�����
q��?��f�JH]�O9��f�����#�8)���'�P5�κ����5��C��V��:�]��zm0���F#$�������*��=��2P�o\���:�X�>�*������:c�?��]?Vd�� ��L��=�YD�~X�dX{�L�������.�G�u�o#�R�RA�m�#܌"�SY���v���zM���B�R��u�O��]s7
i����4���x���24��4"��}��7�]E���g�2"�{�/���Lz�p��'�,A��R�q��P�HDIr�|���B|��T��0[��
�N얝f�H��M(6��i]������=�������nQ�7-F�w�2�ls�xz����&1��ĎZ��pl��p�'�ܻMi��#K��
�͡SZ[I��m�ݿ��%��[�A�}�Ƞ�+� `µ�px]��~?��:��|��td��mKT��L�DT��$o��'�`X��ȭ�����M��:�6�)������pu���4����H�g�2��ҋ��Ў/`fH�|ۯ�`>����B���T���Ac�����({��%�V��<��r
�.D�XOZy �j����r�p3���c�k�%��bVE�ҋ����&�3����E�A�K��}́(ҳ��A;h����O��lqb�v�nH�[)(o��%;�z�[ⅫӰ-�9s�	P���Wk�p�I��Ty�X��ej�v��%��m�9d[�n�X��u�FԔI�ٿʤD`�Fz%��1��x[�
s��!��+�N�֪n{Xowgߩ�K��Pkr�}���2�)2۾�5>�ԝk��;H��[ڭ��su�D�mr��맄;�����L�y}�<Ӆ���ǒ;��2������~��[D;��2��D�I��+�L�o�C�"�b�o�F' �����aY ��v_GW$�|��v�!�j_������G�h3 @����_�1	����~���BX�1Ȇ�t��b)�"��g֥hu�h�)R�3��9���7�#�1�e�(�͐s��DB�YM�n�.5xa<�;��Z��{�=��G�r�a&�����Ĺ�F��C��Dة�y�L�^Q/�G�Z$v�y\����@�G�O����.����q5Vc�K����p��:~�6�گm�ݎ�8��l����z�K�AH�Ҋ=�$�ݟ^uM����:&�EGޘ��*��*,�|��rUt#+|	X1�:B,-)k�{!��c����u�j�m����t�f���&*�?��_p(�����,E����D��M
=���'̩L���� T#��}jn�������Ђyl��J`�hs4�ԇ�-`�rעT���t̸�h&�;���.���"�B����
��)�b��2�<�`m����Q.�{ў�;ȋ>t	8' �J#�L^7��p���3ȱ���^��CTF>N?Į�Kd��i�ڛ�Ɠ`ǖ�'D�7k^���w��
Q���AT�y�|�FA�:�t��^n��w>I��fda]�<%<�z�R��2��9��0�3����D6�0���x" �yH��o��؁��ɴ��娿�6����$=Ypr�Xr��Y���V���1�7�1WH�/�)���Պ`�_�Y�a�l����^�ӎ���y���%��s�t�g|u]4 G���}\}�P���c �r&y�F\F�^,�a�_�T��|�m���!���|4	4�����L�A���"�m��̌`ş(3X"���,�8��鼾�� ~Gw�I�:;�������x�̱YJ�2ڄ������F���s_� mQ���T�x�}%
Z����:�q����:6ި�Ӱ��~T�_�����|�!�xMᵿ~j�G�QvG�@��ܣ{Iڽ��ːUJ�07����'����s?��m8-q&�4y�l8_c9��� ?�j��3&]�_��S`q�5ic���{ɹ�C7[��T{��d3��J^�#E�Z[;$�<�'�SCst	���OsVR-G��
��e0��.,.�~]��&hW��R��0Ѧ���C�_�G��F,-a�4k���]�����oʙ�vz�Jn���źLX�F��13����E��Rip��%ь���Y�4[�y�	аH��ra�$Kj�]��.�]xfd@��P��*[%����ʩ�Ǖ(��Cl��)��tK��_�|�a^.5����T�iM!����S�-�덽@�D,��nx	U)��	: G��:k�u��h�ǥ�ʀ��,�.�㞸<� �2�p�(��df˫��A����װ,��,�M�ix��Fw����rP��ψ��֥����Q����$������r��2�;KR�C����:�_dM�G�ZBNft~��X�״�j�O8$Ǉ{N�iS�"7�֭�GArx�N�n���7&4Kp�8�̥�.���ʃw������ӓ�	p����
EY~��e�>.�eEK�qFP��
PfP�ؔ�/�H{"f�2^#���x)��1��|���Ծ����_�O����[`	�P����6��I`iFޡ9���%�A���*�ݚ4�Fy�����hsE���vM�8d���+xC��n��,�Lˆ$\���F��C.�)s0=)=�'��mizu ���0K�^i�?�nv����w��99�%�npG�`���}� r��a�