XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7�8��,�G���\�Ln�Ή�<���)���0X�� �����f�!�R0����@�"�}uEȮ����3�w� �?�}�:Kj]�Dn�(���%��.{r�Y��op����5fÄ�(��-�m�ڳK�}W(/�K�A�0����ǅs
�Z#K�QגO�R>�&yޕ�T����8՚�Ӛ`d7���v0�X!��%��W�Vm���K]#k¶e:
�������G!�D\�9q��� 4��ډ�j_7^�����Kvŕ7a��[��$rvw+P�cE� w��
��|��䠖*�4⇿�UL��$*���
�H8h�a�$����FV��cE&23eCT�*�*���!GD�p"���7(�7h�ɳu�^�*���kޑ0ӵ+�z(֘���	/���ď�/��	�J��M�O��t��)�~=�	�u�[�=V��#�3��t/Ԫ��~됚z򴋥/M��Ab�Ci��}�x�n����a�CN>�;� �����I%CW�5z��=��`̺@�XHk�!��\�V�t[ұ�՟�0ZC� &L9:����=���0��y�ٺ;���caߩ!���0n^��b/v^׬�&R_Hu���MU+Y��0х�R�Ԟ2�3�gP��U���������L�rY����ӌ�r�mӠ�,`��f?PM�;���:}�L��5�����`����Z��/���ܷH�)0�z6�ԝ�UY�L�s������y(�W��0wt�3�XlxVHYEB    2f50     be0�4�j���j.!�!��*g_ƣ����N*4��	a[1൲:z��y5b�DE}h�?}m6�o��EGl.K����&��O�W~���ED�:s�ï?L�͔A���q��x~L���4�ޒw�?t����@u�BY2-��)����g�i�N�l�m���$3``�}�{0�EԎ,��C�&mE�3�?�~?J���*l(��:`������!h����Gh�'�h��qGK]�����>֔9;��H���?uH��O�H�Wtc&j-�d���ɐd|2�C���j	F>�:����j�f�[�q�A��t���RE��M�����6
�;J�oV)��TV�O)Q�?�R'�� ��B�=�aUI�t������P��Y5'�C���ު7����'�]����҃��p7#~wt��}d�����M�L�ZN��D`���Y�+byw\�}\"B�3��o��6�{���)�r1��SG���2��A<������e�%_W.�R8��h����\��M��?O㴓0�j�C5D�\��,_��L�8�;u��;�r��q	�,�V��u���uY�5[�b����Ġ��6~�|�V�Ϩj��:��q��8�P��Ja$�V�kM���h�0���<[����x!>fe[�����}_�j��*1:�Z"���\�_.��a�B���.�!/�)Nm�-�:�Z-����q�ಋZ�'D����IQ��/��U��@H|;�I�9,+�8)�EΌ��t�c��V�xO�Y��Ǯַ;�L|����qO�TFq@���G�˭ �s&���E�˚(����bä����.�;����4q�}�9U9����E\�$��1ˎ���j������N�n|d���T�6��ه�j�P]�L ��X`zO#q��i��w>A�ы��ޫ![�k���TM���&#�����<y�F\�}=��?��	��X�ܹ:��\XB�I��|�γy<�6������h�,|o3h��qYP��Q �.6��d����}��yBȵ-(w2HO��M�k�z�V�Nmp�g�!�_'!�V�ț�LP��o �#+�D "y0�oo�&���(:ɍM��+K�E��3��y�|ϲҋ;�́ez�2?�Ѷ�_��Hi�ÕQ��'�0�&g"#�ŵ*Pߕ���,��o$�����6�`��Ӊ�q~I����-�ޔ߶���:�D�S�$9{ ��j&o7Y�e�[��S�������Qr7�jZ�o�*c(@����߁��8g��3iѼ�-c
���H�4�V*�p�Pj꧉���� h� ��sOz��"z�q �a��j��� ���	;�^�d�V�7��3�413�P�(�;rD�%�c]��~���U辠�dd��n����h�Vn�wA����s=�3�<��@d�dy߬
,H�
�C����ɣ�x������쁅G�����9]���f��]�&YӞw��B��y��OBi��χ�,BY&��]�+�Y���p�L>����p^������`|�^o��5�
���b�����gPK�j�π�)x/��s�%l��X�5^^,%�W���k[*B�B�d���4]��D�qm��E�����9pP�v�b�`�����F�F��@��7lAj��ā׊/�?8g���������l�\i��S��| �g�TfI�$�έ�Mp��Ѕվ�G��=u>��O��G1ί��8���l�z@�"J8S����Jq�F�
L�C��)�u�,I�`u~�2$~��t��1`����N���� N-�hz��~Vc�5/f�yq���TO]X_� Ԙ�w�1��n:���.^��s�{l���	���˦5\߆(��w��,<�8.UAF��?,RA�\�g��6��6;�b��G�qZ.+zt���;X�񻔸�ZJ��Ȅ���3�@�k���J���;��J.	��r���U,�Q�?�{�np����c�,�6�/��������+=\ז���t�8���WB�7��8��-l0���af�G�_Q�3)r|�{U-�*Y��hq���`�=���Hn�%B#�W�s���a�uK�엵��r�s�U!Mb��8)*Y�S�$���ŵk��4=\�)z��Ko��1��lCΈt�|;6oq��KV�R��,-�-��!

��]V���9X�ơGy���b�[�Z{
��������e%旜��K����b8��,���1v�
 ���ɟ�C���ck"�01c�ޭ[pj�]�i�z�T2�����!��2b��Z����.n�u�p'���̄�05�4�G;�l�h���.��Vm*;q�ݥ�4�o�5�	�{����:h~�����:�=E�Go'�Bh������8J��Z���*�P��=�] lG�� �7駪$6�QW ��?O^����JzVS�,zo�d���_��첹�[��j{�����nE�N�ӷ�e"�딁��L̯rr��y��Mߍ�K���w�Q�w��P|�R�_@������Q�:�)ۻ%�2�R�(J!�D��KY͘}��O�����	%m�L_�%.޷R]�2�U �<��t���� �ׇ�k�'Y����d��P2/��젥��$(M��3�	�a�x��.-�ӭ�a����0�*	D����)O���8�N���'�=�6�	ڛkX'^��o���Kg-���,B�h��J�^q�Y�����ֻ�Rr�]c4�t-G���V�$td��;�)@Bī�A*r���3�C��r���
�qm�o��*�F�)�M�}M��+�}]���!`�Y(��!�"r¿#���T:��;��U`N3�g��7\�3?kV¸Z���8�[D�K�苠�.g�,��� (ݦcv�~�Z�3����<�.�B΍�ۂT��疞��M	~�r(5j�g�;~� �{o`��p/�X��񳈄��w��!F�ϧ��+��Z�����~͉(��5APd�