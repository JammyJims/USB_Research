XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����@��8߆�yH��-����p"��Ć�Y�@j/N�a���͸�صD��5jV�:��:���P�
�J���v4��Ά�U(懻P�)Œ1�Lq`�:�RE-��͛�I<�ØB��˼��ȘW��'�U����/��/~`�������e�\C�k��n�A����Zq{�e��B��`P�V��]���)�A���H�_SG�0��ks��Y�k�2L�t�XҎ�%!��<�P�꼚]�Z�>�o)�H��N�Zk�:�j;*�,����x�y'ǉ���`䤓'-�Sбg�^��>��y�����3�u/�fz��ns�?_���Gb��,��'��+��Bb\*��W[� �I�tȺ����|ú$�"���D_���;ru'nP��GES�"rR��\���ݥ3i
�WGY�	AY�W'`!-����7���x7�v�pM)&ed���ȯMM�OSo�� ���'�z����xYy��{n�;'��ئ�����CoD`ַJ"q�����KL'�[�H���>'�amO��1<������eh����߰N�?�dκsb�{L��Y����B�U�f��f�k�AO�k�.�qȱFzG���ǵ[id ��ؔ=\��$���u�kL�8�2� W)Nn]�'�l8U����Ӓ/��aZi�Ll�{�X���+���j�%abİ���_=.�!�`0"��Q����~Aۯ}[u~R �.�%T�n��e�"tձ��V�ΞXlxVHYEB    6f05    16703��'wLg�u�a������FP�w;�I�$.K��U�؅�3$�hSS}p�=u�T<8�����R�d��m���H�[�k����k&��d)]��+.�DM©̕с��d�`�wG��S�A����\ �L��c�Cl���$���G�չ�ǅ������ ��FҸC���o|�j��_�"Y���a�sʱ�C�P�[$��A�z�u�� ���Q���1��S�QԳ��O�<�~��}Wm#�����x,�z� ��q[����� ��w��~�uD���� ���n�z��"����ڕJ�w+�^2'��q�;��}�c��@��^��;�����c��΀�R�9�CE~">
g��26sa1�LR�p`�S3���.M�*��5��n�jd�3��)���;�	�K��ϣ>n"8�]]A�o�3�Y�&o�/��5X�]S��˷��]�l��<�n��u�-��m����E	7Ve������>���WI#��/t��:�L*���K3�!�X�1��
�#�䄔�\V��{NE2؇�a��k�y/crK�&,^H
�D��p���Y��z����{���O�����Q��6dHD����3V�'�sP��D��ӻ3����v�r *G��2F���T��"S#�S^`죒���k��������^X��C+2:T��D���KM�_s�h�����*���V��Y�ꫬ�Zt$Ԟs
�8g4�]V����>,z߫1}���ެs�2Y���_�`�7!��F9kv�1=q��4Վ�8�����B�Ò�,j�%�`��I"�'?��G10��>�rr�^�����( �V�6��"����q����iG�Cq�e�F�Ek��{��*܈�����D츦v�S����.�+����y)�}J�Ҽ��EF�iH�F����lk��B��z�eݟ�GHLn�D�����)��1q��S����K�lDl|埩�Z�7��Dv%w�7G�fs둨+�P��̑>�8�*WƖl��Nq�4�_�A�nJ*U�����6"���iX��͟��L�l���^#�+t����=��@U�N�^fn`H��.����r��͞>b��=���u��y�_b~���4�*!I���m�N�+IJ��d�>���?�[S�ϧ�,��FN�8tHz�#g�Mm�����:u�>9��/��E�t�ǧ���*9U�g?;�q��DQ"�!�<#y�毕\m�&��jY�Ħ����l&��u�k6����3#���vҶ-�.�],�+�5�l+L���8_,���}�`�\�^�\%
K:�|��u�:�/���;^�|�9QRHSN7l�y��I{	O�4�)�Z,�u6��fl��*J:�I�ي�ݕ����;
i�2G�U�g����>Y��x]<�סּ�%�f�L�q�8��o�L"Ϭ�Q�!SВ4+��KϓR��'hz/-4���ԥ�oe�!Kl ��T�����d���O�丠��tTmV0>�Eͦ!h4d�y�������r[Q�`q�_f���A$֔"���ХP��fn;!��G�7A�=�4H�!4���"��g���$��ʈ1�����5,���?��8�!�!�<t)�PԺ�WDs�k�~$OI��𬖩_T��JgK� �X<H�:ƈS�m.�윛����u?l�%`eһ����M;m�DK�����h"��Ą!L"�hgZ��-��m����3���X��d�<�o��.ڠ�1��
]���sb�t��d�؅�1�1K���_4�R��G3� ���d���z�`ܹ���fQq�����C� r�C��+��z�r���@�V0m��١̕���	.�c\6|A`�f4/�.j������Pvv+����9�#�9|�S+��o����r���u��&)���-�]ߦ���`~<c�6z(6M� :!>���$f�"0�~�u��l�n�i�=
�������5Z�T��*�m���=C��� ���%_�]on'��,m"K|r��Pt 9'��บ銩\�:Ƈ��w�$׷�͢�ߙ��#>�/� @x�%=���^��y  ��������@TO.^�q��2��$`� A
�2 ��L�I����=�6��%%�s!����0$����=;�~y81)��x�9��p�kLȭ�CLmT+�K�Ǣ��$����zy���"-6��6h�1mE���d�"���/�@��+�aO��&�X�k��$�4>�eḹ�G �o+�mqiSN��^��=8j�,1�n�Oч%˼�a��(�OL3��P�Z2
.͋�M T؇�5�Yq]'-5��vkB,w9�K(�S��N��|��U2e�B�DԐJ6�n_�9hfȝ�Y5hҺ���v�_��v�u�[�tú��U�'�(9C�R�⣡VR�a��0
t;o>��i( 9>���Zn�l����Ϝ�f�!DNM��l� 9�^���2r�Y��ft�B-�Md'�a2�u:R�WS���@���-bx��(Q��}�!�R��(Y�i4	^�!�՞��(4.M������^�"�h���E�~w���L;����s�F��q�����~�����pR~l!��;�N��/^�P�a�P!'\���������	�Z����K���2��W�:�\~���E#����'�r�:�-� ��B��i�H|���'���%�#�@�Ց�m�l�r�/y��1U=�dћ�VnV�l2Cv;�<Yr�f��l=P*7x�ko�W��d��a��xX������uF��~����η	H�<5&��%��1�ث۫�W/�I7����l=JH��xAI1k�m� շɫ6��@�������yE�xļ�}�Ye�1��ex�)!��]�� v�����<�j$7X�ȨtCO2:�m��At�q���z���)����Iv1l�t��c�g��1��б8FQ��\���M%b�#��\��x8\��w�T6Aԍ-���1GajC)�j����gf���.����U�B#s
���{;P��&�t�?�܃�J�f�/
Kiْ��\L����\V�4E���^��{�(���*��PwaYBѬȆm�4DW����6����3�F�1��^�_c�0L-��J����*�Ȋ*d~��;���)�ģ��d���f6�JI�q�v�.;������J�1�2�fK����C�$Ά�����O3{G�f���m�Z��V?`*��1�A�X�"��ǀQ���u^%���'��1)��C�SFԸ"��]�B�����O�=��j�f٩z���dC��8�=C��;N����H��q��D��V�V�(j9�|��=ǜ/�{-�1}�1Z�?K@�޼����-����n]�Ii��#�tp�Kzdq�Ol�X �� ����0bz���k`���c�)�ea�!�%���P+�=������2�[|�.U��r���C�G�u�/IAP��Gl�q@�f-r�n��YJ�bK1����J��.C��\��?�h�� ��|�T��3��iR�%�v�3n��Gctr�!9XS��[>7����
!���sZ��FbZ6�vU�9�>o�菹�m�v#�=$��� ��΋ME}��Ux(|>F�0�yS��P�{�K�V�]������2�H�گ|����.À�qZ/�Sb��p<QP.p���0T�C��4��K������7�H��\E��&xj�'*BƟRJܧ}�����b��	���![�]ʻi��ɲa�N.O/�7��uJ3n��)��l'��f�{�>�MV㏓A���96 ��X�f�&�u`�`gWm�t�� ��,����Lhy�3��>�*9����(o$�%��d���&��q�Y%��+�9U��z��y���/�����9�!BJ��V�}l	���l�6Xr�[0@�&�� @���뛡�<��ς��8j�>r��'$߲u� �!���οjp��B�Qn���mҊBq7��}�����l�ԕ�]�v�>����^�W�6��Ǔ�K�o�K	���������!L��2j��d�.}���c�2Rޤ�xfjn�7�S�H�jpՀ����m���V"�T�)��̉�H���ל�El4�*L��e��䫎��r�R\<�KqP��h��;5��{���w��ț�6��5�����r��p����vD��|�����;����K��R'�1oM��I��Y�ô�ӻ3�V��I-f<m��i�z+͜wH*5+i�D�����b��8K�Y��ŃE:X��,e�����TXd�)�a�l���_,+x�`��{m/3b�s�ň�sj��N�i�)亀�Ūd�;��[�v�����e�]V,c%�0vސ�g����|0}�)����$x:����<�2%�$�֎��ij>
��/��� �U{J��9��{�葚�˝ژak��0�����vA?&�x������)U)��H���x�
�'k���pM>�Aqe�6�뗊�[�σpi�_���7�p�k�C�(����F�M
���'w� ��d� `L��g/�*u�WkX�	��Y�� �J1s��`�ͣ����n���%�HIZQVJ���!���RB���G3^;t#0)��䡦1���l,�R]"º������k�P@������H��Z��k@����I�ƈE�]x�H�u��Ȇ��YE7�(Qi*�G� �k�7]��v��������#z�m��=����"V��B�%��pd��?����^ݧ+:���M>y�y��*"H.H�r��N9��>sH<��h.��I�G�%��M��tlP4A�y�͸��s޻.��d@?�7�j��Y��P�-���eQ9j�n��̓ ���w������7?�!��;ऺ�Q����M�(lSޱ�=�}���[+�uwp���2Ƴ��ihY��WP��LF�D��z�o��P��	@<|9*i��(�����(r�ч.Ҫ����>W���0K1e-S�\_�=�O���P�"�Wq�d2af��e�<��aB.��y����V܂����!o5T��Ț��S��yu6%B_m*�O���y����;5��7e3KZQE}���P��[�I�r���Xް���mi4|�A)q2�⹠${t6���,���4Za�~�Į�b1fh""&�.M=m����B�*�&�Ъ�f� �j��|fRr�k�-�ܨY�3i�r��v&����5�3[�!J�e>��o�+e=�Д��H�.��|���JM�e�z~|r�9�CvCK������R�l�l0�����3��ݸv�N�5�~����΂}�o�C��z@�T�c`"2�20n�2��L���>Q<�y�6�N�|�p^�2�3=��C��vT��ם�$)��\�@#��S;P���L��ta`�-��Q9�<�(��J* j�"<g9��c\e��T�'�<8Uc?{&7�Oh
Y�l�%�M�8����Do��[5		dZVlބ`�� v^��ɳ�^���{���B�>I���S���v��dJU�+�g��{ՂdW��Y��:D�(0Y���q�%�#���Lc@t!Ұ�˹�:�7� ��_7�b0}31]2G���Q
7#W,貯٘�޹ ���dO