XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����.gמ��GE@����A�s��^�?͈f] ,t�a�lo��%7�ӥ4��ϼu*~Z��fʅ�n�WL���=iQj��u��4��@h��`�lS`6����E���yC���:���¹�G�M��ji
���%ʵm�(�/s4�rʜ�u�c�B������]�5�"����Co�t�u���yE��l�O��Mm�(�����+�F$���)�,x���Z��|�AQ��	�z��$�����
�NI1���"��23��Wd���� `�dB�O��b�� �
�ڔ�pN<�WvhoQ�z�`$�k�"4ض	�
�v��v@�&�+ID,TO�d'R�c�.�C��N j�h��H�DC�+�Kv��m��BM���T������a��$�>�%ƻ�E���~Z���������s΄�5p�S�N����5la��)���7�{(T�����gd QC���H�����+p��>}w#u����E���P:#W�@|�g-b3a�R����BG�BTi������i���߆���9@G��NXKTfl8�>MX�@�,v��rF��KX�J%{�!�S�X��}u�fQ������t0N0�y��Z��Yk�*��5h��KФ�C9�	p�_��d�Է����J��
5X�D�^?�;_�3���h��!�aySG<nNF_���ˈ����~��62�����~W��6ǿ���Ӻ��KJ?�sJ��Ŀ�V�T�[��f��کNt\�t���N<b�XlxVHYEB    2bea     d90g���+]%k�3d���Aݴ�'4D����A�_�>�Pf�٦�fk^�[��{�Zlc�z �z�63�I9Q{�be���G�l>]�=�ؤT�Ȗ�r�VXҸD �"F�ҷ�-Kwn��С��J�kV-*��o��vy���i0�����I7�~0�?�`|�����c)0阸�Q�:x�eރ��p���GV����� eUș���c|��<9#F�uƃCQO!bD�{h<������R�S����n�?˸��;�Aѐ���-Ǻ��4�iӳ�����H�=XM���S�՛�2�~^��v߉-L�^`�o!�!T���S��MM�9a�N`gҫN�n�?f��W�Y��o+eDC&*�L�6�t��&1�?�Λ7D��-��>�V�N�����4W3Ԙ�5�j�Xd�	�`�,���.��x8��]q��-�DjAX�@��v�e�W j�b�hlo^j�V�{aW_0d-��vTz$�G��BS��BHA��>�Dd덱�u��+��1
���9����p�O?�L�.��Sy�\N�_ԃR�(s<���ݝ�r��b�!�B��� _��o����Q��@Cș﷽-L$5]��	�j�˒%R�{;�#8��u�ܠ�d���e��Jq�\��uk��5������n�.k�#:qgc�N�.:�$���~�~��6R8J��[�.�p�-H���=w��U]E�5� �V�+&<�h=OP-����>�Q2zu���v�j�c�?�?�t�7s��� �9�P���jZ�A&B���M�#,��1�`0�O-�P.�e��0z����^=T:�J50�f ���iu���.���!]+f�L���6]�����W�-�C�b-Ih���°!�`ā}�-9T�AGX>>dN�>6���HЧ�WΣ��N~�m�lI�f���C���ւ(��C���F�6_�p�+�
jݶ/������9������A�����Tu�p�&k1�Pi�!L�>y�谵�=�M�q���[h���f!����]1��7�a$xFo���� ��(�z}�V�H<m���a8��y��~�k�5sJd����}��mxD0c�n��FTb0lʂ�u@���ȩ3q(�6��/�0�L���1���&�Z��aى�4�k=82!��r��g��*/� ����t	`�h�*��r|��c�t�J)ʸ�vV���G���k�#��ճWN7û�(v*����'9Q�%�ɀ�ua��cc[�/�l>������$�2��,�(�c�|VM�2�����V�R�)t��-M�tX��mpe��%iW]��2C5�ʐ�*���[�@)�Q_�R /�~C�P�Ԩ�o�*�s;�T�������6
�X*\c�s���T�҆�t���F�7@���^��%�`J+#�f��7�0�kQ�I�_$*�˱�>@ 3ڦTO���!1�k#���-��|���8�>Qq:��[��p[ΓYs�C�A���8�̤^<ar�P�R�����Vf���Vv��*���_�qev�;����(���◷\�H�>��(7��z:��W��܈�(��f�~/�O O�����Q��+ɐK�@���� r�d$Ad���bùK�,%
[w��]x��#h>��d�%�,����U��5e�X?�m�v �CeJ��Z��4���p�����i)�判Y�߶F�B���G�b\=�F-?�̂��н_���z\֓�v�Ci!�Ƀ���O'Rۥ;�gaG�S�,E5�Y��'=�Y���N��ŖHA�EI-���(f�iG���ֆ�����y��R'�풲?���g�P<��h
6C���kY�vL��Udx�=��&8����R��VP[鮺ɬ:�ެ�Pc�5ƫl��}߉���_YB�sߙ\^�J=��
��� BA���⵻�k�e{,z��r1o��Ug2k7��6G\"��T��ۄ�q"�����pb��͋����,��Wv��|�r�����������^��
���y�Fm˶P�`��BV<���-!���W��Q(@t@@��vs��B���1����~�� �����������r�!#�9��|�*�f�k����)!nTFQ��(8|Gk����P������Y@���>՞����y��Ŵnc^�i��Y�EN���{�����a�⇲��i/`�6�ZhV�F5h6��4��c��^3;�	/�c��N2�A筘�9��`X�<�R�C�϶ϴ�,`d�G�
�2���|��q�Ϧ�Z��W�&���؂=��y�HͭT�(��J��ow��. �MӶs ��?�9]{����kᅳN�c	�=4[ao4%��S���������տto���Ő�*�tv+u��Z�F�x�
�3�������7;����?�1 �^%���Qk2���K7�]�e:�zM����~p�����XF$5@�"�^p�A3%��o �(���	ZY��8�����������H��7VB)���p���T���/�@%���"�5�t ��H�E�G܍m�W	�p�����J��I�]�] �˛�	n�S~��[��N���tkpZ �Y�.P�5�k���#g1���7��&�
 D[,ɳ�ҳ���7�5�Z!��.,�u�?*�>�D��Ur`&��A�!Ҹ�1W�*떭�M���hm�~9�ݲ�܆qځ�O4�����ȩ�@ �XW1zr��R⻊����e��X�B@G�P1��b�ظ ��ޟ%��p~�\�:C�2�s�z�a��ؼ�Zו����x�8��ۣ'��P��It��:�'�9�O5�ا�
��e�ͼ��u� �^��d�po���-�8�������a����5��I�����0�y7��?t�T��\�O����I���;*�^��̲��8�B�=tt��'��2�ؐ�C���Z��-੓
�4>.�(�4�<ݟ��З�hU$}TP%-\�����7գ�s�s��Q5R�MF��l&D-kG=�S�0�W5U=-��#_ 6�x&�-͚�<��J��Q� ]Po����P��Ā�!G>�����w����gL���W����!��W,X���߅��LH��zɤ���E�>���~���_"�۝[}��T+mݰ ����I �T=���1hMǃ�{����[@�z_��^�a~p�4h��u�ҿl6@�fyv�pZY�\�Gx�?n��R:�����nF~[�2*��=�	��{��c�Ι*4~,����К�$��Y�қ�k��VVx ��k����dsg�-g�͂�A�� �'i�E�xS���{�t�Fa�V6�
�s�����Z�R7��B����je��g�mӾ,�e�3��Fm:�����z��{qt��H�2G��dlW��6�yH���L�؎Ã[�����e��
