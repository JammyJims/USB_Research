XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'t������c�bl b��TM1�{��.�8D�C�L�J����G$8�-9��Ώ|��6
ƢW��7v�ir>Et:��i�:��L:_��BP��ꫠ�4
�)�/�(Z�r���*&z#�D���"���N�X�x�@�x��C�;q�����d�)<�Y�]��g�Q��=W,l�[���0�+۷��D�0��j��Ͽ��n�9�KJNE�%��^4�w���c55Ꜫ����Ɣ�[��lN��;\�ۇ�b���9���Uuȧ�zq�V�����^$_����P��>Xx�▥,Ri���WЮ��4��by\"`T��R�C
�Z�Vo���B�[��)�ՅX
v-�ū�F�'������}�.V��چy�phd���G�6��W�̞/m�z��p<54�Ϫ��A>�
gh��]^��.�ޣ	�J&e�b��!��r��s	t0ۘ4���DyFþ�L*�P�BrC�1|�p%L�l���Հ�}�����`qJ�aO�HFk����ΌC`,�{قe]l�U�a{hU�L����.��0�)o����8�d��蚳ľ^��"�o̶�s�Ϳ��#���Fh���%�u� �p�ӛM�H�+��3��]��w�s�b�)%�sb�z\�~Z��	�pS!���_b^�ŁC�V����u�x��!�U�-��2��bC�s�;K�!�g/�y4��!���7@�����Ńp�߈哦B�x�}��w�G�P̲ Eo-L:N.�/�3ͤO��]ٴ�XlxVHYEB    51be    13c08Z+� ��3�<o�����T(]�j���(�.��sZ��79N$k~��-$�!��˦��̒r@k�U �}Su�r��?5IQ���e�-_\+�}w�^����z5����3q~��!���"�������a�&uq��j,2(����x�1w�Lh�?0���J�Rg�T�80t�ê67	��D��\�q
*��l�F��IU��l�V�@T���!���������vC5nZ������?҅#����o$���W�4�ݙ�=��fк��%�=�v�����C��9#�t�t��ȝ�r��̭��e��L4R�"�R}�J��=��X:M����1e���u��! ���_��=�ks�D��Lk���EF0n[|ͫ���b�����$/4;{k��-� �«)���hLg�{4qm����vr�ǿ?�`7��3��+2T?�G��9�n���&8)�ٻX���g��o&��S��R�8c�B�`��\�k_��=���>2�R,N�`�w�w��p���+.J��ݟ*	6#{�Gf�xȢ[Ш�M5gɞA�Qyҁ�3�6��<l��k}@�ݵ�r�w꬀��%�'�µ=�� ��h�R���;#�e��b��n9�D����t��f^#�q���e��r�~��D릔!�Bt�;�0'�|ő�F���n�9��,��o�L���&�E��AiϺ�¿	"!{���Ek��o�Sʝ�����K�>� ;DO�vK�q�K2YH/���F��n����uɤ\\�}�*vO�)o'�w���#�{.�w����'�-�	�2T��xч$b��l�!A���ʙ�߳X�t�9,��7:��'�����d내�Wk�E����(��i`Rւ������>�*Sdʕ��#��O��R�v��"e�"��c�V
rM�E��5*$� ь�Y���[�D��W&�k�Ę)>��O&��o$��*��@��R�r�L���Z<�����N����]�:��1��#������Ō�wƩv/H����'�}��tL!��ʅQB��r�í�����F�O������N��L�G"�	uo��(E��=� ���$��4Ym����P�{'mE�YB���T����#K+�77��B�4���T��	��fW˪t`ʕ��D��,b��w0�)Q�QU��]%�g�A�k�@��S8{b�_�V�F�����Y�g��w�ի�f�t`ni����|�x%JN4��� �]յ���ի?h�TŶ�2��{�XU�.0p�������|�䗮]"�)�:�.r�є:���գ�Q'��z��+���V�Q���qd�z�������~������3 @�\����᪞�O�˙�¯	-q�t�g�҄��ʵ�un�g�j[-�;���M�W�tԒ��D�8	�H�;g(�I�7c��6�"�c�VyI��[��J>����ú�
\\g��] @�^�j󗲠ˌ�Y�����
{���I�H��4��cb%�3 �?s(&�ݔ�E��T�LuC���;̤�9l?�����g�F�6l�����h %�@'�h/R�rT����&��_�� k8�V'���KYO��QLA��Q���M�'2�=W�"Ks�[F$����P��Q�M��	��T�i�ȍ�x�&��.�<�&�T]�W�s&����v|����n��Č�ѧ��
G� C/�� Z�@�5�����$S�b�튯6�Uq;�ߠ�F� B,��ݙ��m�~���=�n	&��m�wl3�v��y�o&J�/��>wڕr����;�P���<-h�����m�G�`FX�-@r�P�:%vl�yGh���%	P�bp��bYh�}��`+���p_j�B�J�"LЌEO&����U�����tL���N۵:���V�>���_$�sf�zL�Z����1'u5x̂��S����V�s�Ж@f�����sV���s�����et�bA
��y�ʲ�)�7[)8�F�J�ϲh����̣�A$�,�b'e�1�ڪuR �3ۓ�l0�Mƾoo��>L��R"� $��I�$ԕ�a���on?����|&�!-�,�;��y�^�r�QfVL~�|Ԫ��2pV�4J	����sܙ~K���Y*q�+���K
ε���ʽ�K�8H��>�P��,�ڴv�������3B��e�\mk��p��n-*����2MS��m�2�L ��~��I�,��t;��=!�'�L%E�T�����W�
���h�$߁Zk��˃�ڔ��y�;!e7��nP�7s�:�0�
{��x�,5[:mZ�`���h�㠳c0�u�����6N.} �d�\c^���cZы�g.x��t�pJ�)FjSC[=I���]K2���yP�ڏu>緝1S^��غ�~͠v���y�Lwq��=���kYcUqc�����׬��v� ّ\��G�R�o�3g*�ZFPɁ�ԡ~�&���7���v�{���_J2�:������f��y�YN�̻�G,h<ƅL�����Y�-{��^�:�E��	vA+���Kiw�r�h�j=��%���M?^�v�<��xN#gAp~2GB��dm:�פ�:چ�?���4�8��5�?�����P%�)�,>��tKl�+3�vt3$��ga�ښ�{H�4�C����GM߃b�S���|l�-v�+Y���;����R}l�Cݴb�L-T���5a�r.������*:��1(ci-�-��9	����;�!\=�o��SE����|�8�Q�Mn]Tn;ƺ*�S`�ڒ�6k��;�K�&gE ���@!}�]_�I���߶��v�L!=�_?�5��Lnf��ߓ����0�5#��ߵf�h��6i�++u�cf��Ax�J���4�cZ�%_޲�y�CeΗ!����Tȥ#M$/e�G�w���$m�/(W0�,�(Ry$�?*���3T�hT.=�`iv��#4�@�������7��w��`��W���-�^h2�x<u/]k������I���pO�\,�����<�<Q��s��@��{��]�]��%��^� �B���ۙ&g6��s���g���`e��|����A]l��h���ߔP���J���-��<[xȲ�,T$�#�{/��̹���o�a����b.�3
;LJ�=��%?
�xb}h'u���5v��/n�,���'���>q��+�|�J-��c��.s^e�}�''��n��~2����y/ui�=�}�_��ٱ��,�fڣ�P����ʄ$F>�<�F�*�@�Wf�?�� ���ˠ��Y���S^��fb�D�EUΠ��R���r*���-��w-����4���Y�����"s3G
B�7F2W��n⡨+*qE餘��B�FCҫ$+}�%��I	���"Ё�pEB���Y�?>�%ǱZ�\�����i:tW�}G}*�UJ�CMZ}�� ���г�I�$ў�	��No���`�֚`
���̟�I}��;�)E��	���Y� ��'��h���e:Z����n��F
â�^:��;��~��ɍ��#LMUOw����ώ#n��/2��e>@"��6HԲhmq�W�Q�N@�'U��7%���Q��O-��k�Y���XҮ�tf�p",�z���� rN,Ԅ	�w��J,�惎b����=k�|��>�ږF4���|�~��{��f��2%���t�-�٥tnS�0���HW��\5x����Q7'�=����e��_�B���f(L��lMsˤN"S7P7v}����x��(������*���Z�j{����,P�!{l��9�79jZ1�����\4��r��Nn�p��k�sޖ�������O�O������w�"��a��k�����b�����xc�
ch)��7�W�-�Ne���R��ܱv��R ����?���8�^�;�KB�:���:��`���.�p�cz�P�N�v�0B�.�9 A�O���i��i�<sw��ӄ������+sV�'���$В�UB����l��Q�g�RG�T���k ����9�"��;��>�H"����om馜e�N%������j��ԙ�/�-i�����b��rs�l���B0����ry������`p�!��,n�����������������(2M��r��d�lN}:���������s镲0{�b.a�F�_����|�%y��)��~(Oe��-�
Ў>�U�0�d�Jh�D�yq�@���ܮ��0弢�[��<#�<�n�욀 #/�:�9�qJw_t����GG��ve��J����_���h��;Ht��匠~�Йv��	V`�ـ^����.Wn�^��T�>��H��e��1]_WL	Q��x��[�s�E��@�H��sRce��;&�B̖V*q�tp�b���Q|��g���%��܉0#ތpw��a|"�m��nfu��1۴�u�eo�d��k�v<o�W�����S�y�5;�%�!/�P��1�+b�;$aܙHHYqd*�%F�z ��ۆ�x�/�'6ȦxC�"�@���4"��>��'[�����يܷ�����J�xt�g݉Q��9�ؙVT��T7N��♩�ס��H&���*c,B ���S� Y]z�xW�S�.�v��lm8_�(h������C�1��
����+ُ�u��90�~���X�0}��+e�D(��e��:��SG���}E�t�Qpj�6K��Lq��Ν_��j�.�b/g�K��zr�3z폽+s��"��aC�2�"�y��5~�����(	���Ǭ�-S���Vt���:�Z�C��{n�T�T.�iSv���9�E�	g�2�^�&I^9&�mm/M�@�x@��$"F�,n(m�����:;�M��'���.��ʜ�>���(����I�]��5O��1(��Ĉ2�H���a�y�f7,�F�ݿ���O��t{aP`E?��քr6���R�k}�v���Y|V7�".#������	d�@��r�