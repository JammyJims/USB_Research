XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���eL�}d��'<�L�(�De6R���f�{a�r�N���R+�.�*��*rT�U��D�]&�Rq�%�jϸ�zlJV�є��/�%io�#gq��`��i�2�z�x:	Q�� �6���^��?��e�.�V��%N�ء_�R�("vfs�,%�ܛa��V�pp6�|�v��|-�s�F�/!f%�W�"q�Ehm��ǅ&F���P ���K�tpG�"&hj�-�*�!�y��o\#��L�t ;�E:�*��ZB�J�f���Xɴ��0�H�I���p�����ȤG�v�T�'���f�Ve?�>N%���Ȝ�q�b�)���/k<B����,���0\-�WG�ɇ�Y�)�e�a�;�L���cW����SˉiYuH���/��?�����:l���inF+�ө��_�.�B�,�54�lX5������ $#�l�<�ɘ��hN`r̾h�
F?�A��9!8l��x8\�S˭�?�X8j'@�p"dq�!����Vx�Nc����`�i�M�wr�*�0�&��.9m7`��{s�W�S�	"�@c%++{o��C�8���\	��p�z=oy�1~�FB-�hYFg����U�/x��2��Ϣ-l�~���������-�-i���lg���WYԉ����WD���9�!�S��f҆�6��%ʕ��ԋ ����T�)O��{�)b�LlR��Ƹ�DH�ޓ�E�|�`3�}+Dz���Y��iI��qL��ܗ��Z����Y�&�溆B˗�SS��c�s_:�ɇ�5w�XlxVHYEB    2252     b70�o�L��R�-T8V�x�5�Vd��d"*K�S�Mv٬)�P"p��:MI��7�n:���>���ƿ������ ng���*F�
�%g����e�������L]�9��%��ɢ8mpɟ)ӅU�1���uw�w#;ɝT!�z���
f��\�m��2O��j2}$Y�R)�4�3�7&��"�@b���Si��)���|�{	��>��ZU����:�7P3:Myc��x(bN��K�D�����gZt���^&rŵXDO���9�jO"Z�Kh	�3�iR@e�s�64Rsۇo���������ZG����������[���]�1�*Sg�����;uE%���(\QƍD��v⦅�M�j��E&`y5�I�Gy��댢Ʃ�f?��J�Bg�����J���M�i�=��\�S��'�m�2��d�ErÚ��]ZѠX[%dN�1!��ZW�s�w�y������_}���B�v8��c�������0�<�,���4!�j>�j<
����7�ĘF���s����=��M�Ђo����*�|��Dٕ�쀜5~���/�$*Z�F��@�Mbr���%2ā\<�ⰷ@��KAmu��(XDf�Yid1T�2�����W]����
9��@\���9�Ě���o���(�w�탵mXpա�|:�8!��M$����M%ҽ���w����'_�z�_��08�p�Ld����8(4ߺ	:u�(�8��ɠ������B�i��!B_��7�Cѣ����k�y���<Ƚv�2��b�w�* K��~�j�hy�Q-��F������~J)1��Z��'l� _����b�W����h��K(B>J�k��e�fM�B�t`PU���rS{��W���8�6��FjE�K>͂פl"�t�J�0�c��[�{���s0�喙j�e�0(���(���V�;B�آ�^�Q��MoJz^��ږ&��Z4�����t2��+,)n�_��Qq� ��b��*�zU{�7����\K��n6�Fա[fUn�]����Ze�W+�p2��^�Y����&�O��5�N-H�q1��{�0�����{롖T�j���-�Ι^���H_���g��x��4��㸈�X�$ߨ8;;g6H��b�$�\d)�v�p�?j}
�*t��a�jbN�q�"<���tiя��Iw)��1p$��{��hOƵ��_`za^���6�+�ͦ��[M:��Y�?��ĝ���{$#��}�K\��������٫u>�"�t��i�
�z���y�Wo/ٛ���ӁƷP�oh��X�6������p�� Gc��  {B,%���GV�gRX4:o��Tm��{��-_�\��֤�:�lS���^<�Ϛ=��g�9HY�qp"��]R("v8/�;�=_F�p
ˍ�����W�Z�1����X}�������*�ŊtK�r0?�+f �^b�P"4)���H����WP����h�>>�7[���ɠe<0ûh9��)��O)�}��0Y��&�3��O-�P�A�Fgۤ�yv�@xT���&H�}���_����n��+��s̤�M���'�M�͠�Q�*�3;�q��[�=��e��V�8ZE[�t
��?��"p�R|[����1�H�Xa^�X�*��(���`ΐ<�F�d�s-��Q|��M"%��9���E�@`ch�<A�f�������k	_·}2�P�f�2z�2V0e���7g�^�a�C<����UE���5V�_��Q0p��^�=
�@�f���`o�Q��@::�����'�A�S���^ʎ���l�ٞp<H���Ţy��W�W�&=�~'4Ydaqrm��^�`�dj�)����a�}��2��.���k��,ZI�
M�t�xs�ܦ������`��v���3�����8|���G�u�R�*��&�S���v���v����L��6�/�?�#��>-Q�$f��;co0S>K3�!���A�[�����PȻ$�I����˲ TR	hy��O����}Ƀ��V)�҈��L��f;5ڹ^�"�N�H����o��۷EM�M$s�ܧɽ�I-p�$��3G%��?1���ᵤ����a���؃°���./A<p���5Z�:;��!�q�]�5��B=��ua�@��
��.�r۩"�!پ��L��G�:��g7los���׍W�o��=O���D���oP��k$S���<iUt�
�{P�s���MBjU�:ӎQ�V�4����a�f��b��(j��WN�N��o ���;K�/���eU[@���$�W�f4������=�-������ˎS��q�z7�rl �?���	:�W�
?�窀5Իx�9��3�h�;k5�`�j�F�S=�n�4�8E3P����a
$��Z��>E�lq���"~�<���ot��4�^X����S#͘&��& 7|�p�u}c)��i��kˎ��R����y���?UK�KG�$��"R�.�6�e��t��=/}�:����c���`_�]���DtJ�5i1��3$�.�o$�� �[����H�}��*Ke��ߓcǄM�B�STa6�7w�oڎM�p�Mu�s�qy��Z~=4H�4�"':��8�B�t��^ �g�9�.zyu��e�~��������-0�����0�iXx#�I�YG�3Z˵L�qJV4�@4/����N� ��p5�a�ӊ=�u�x��č�u"Σ��*�8M�����9�i	] k;V?\,���׆<A��Q:QF��/)�+�|녕��v��t��ݡ�6��2S�!�Jٍ	��!��S#\[�-Qv����� ��f��[h�I�p���	zU�{���3�kt����E^P�a2���x�M΄�H