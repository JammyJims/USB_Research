XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W<�4�r4<�<�^������n'�!nm�qnG��͐7&��>*��K[ɥ+i���:FI�4uJ�U]$�H}��煑�~?&��Z��լ|#�hQA�ҀB�OO�Y��,,tI7����:4�@�4�+�M� �{S$s��)�f�\~L*�}:82��f+*=W�E��k�LaF�ctߴ�D�`م�y+"c0�	����Ne�y�b��z��=��z�C/� r��(>��#Ukip���xk�ƍH���(23^�.��>.aK�vF�ގ�*�4�Y'M���j������f0' �7�	�tv�P">2DpKzRZ��OR�jN��R����h`�R��pN@���I���y9앆TMXgTP�!цՌ<��g��7jHRV�t:��_�j��$ߦC9��V&��~�K^sW0���ؖISHo�)fc�X�C6�W��f��)^�#�P�m�3��`�>+K�C�g�!r9�N�+��ܩ��h?݄N�1C�m�5�$�WZ�R=r����B�%�ה-i5#�02��{�W��HM`ۼ�<���x���x�N#G ����0<\Z�}��W��j�H���;�U;j	�>�I����WA#|��:̐�/��!;F��g�pf_��"��k��F���_��D>�U�a!|;�����C�S�8��A���	�\��cH,G%�_vUd���:��� V�W`�4){�������zuoU��no�X�ph�.�Sk���j�O��Z,�*���XlxVHYEB    58fe    1550�/�Dz(�o2��[�ہ_���9�盷`�mo�G��A�j)􅳉5E����CC���g)���~%��{�߮���j?('�)��Z/��O������d�}�L�J;�!���X�j:�ԊS��n�"i�A�hEfu
2�d� ��XD��T R�D\�J��IC��4g��M�o�rlY 5�����i5�F*L��󅒔'g4��iǾڀ�����W[�.�R��׹�J�Qrw�j��ܤ��މ��.)Ѥ;N��7�@.>����,��� Q�MlL�t��W��ρ��a��|YM�B���DWPwHY'�t�~ʿ�������P���^�6�����-!E0SӞ��K(��X@���"�J�Y�(b<�y:��*Έ��P�  (��,�5�v��-z��kc۟H̬Ky�S�r�PM�ҤՂ�סF��t" �򞱃]樒Qhٵ�uת��|8O��$aʀXa�nd
�S�>ƅz���0���~�2�LW�]#�i]���ZE<~��1�^�c��W�To���~�ʝm����P�x��E	)uD=ی4i��L�7Mև%v�*~���۬M�8�����8}���N��s\��sU�y�����me��'xn�[�����T�*�c�sDD��P�Ǳ��p�)IZ+g�D��W�Ε����6�d���:R�=���ܐ7��KE���� BүL�h/	m��,���\�	IO���?����p���H.;��B �*oGSzD����)�Bķq�:�4#͘��m��T:�h�Xᤒշ]��ʅ�j$��<��DZ���c�'?y��^��GBET|��!�qql��"���r�����9)�Q�gǠ�5я:"���%�Ϲ/���()_.�鞳����h.Su/ftbN��0:o�i�p�� 	�RG1���po?,�We�B�Yw��d�bZ
���OnW����ۛ���T� 6�n�Zi����F����v!wA#�;��+pb;狊/���n�o2�S�A%���i�ި1R�������d9���MJ��!��$�}(��jbn KXgL�*����T�yGߊ��"u�T���K��eO/��gKS�D���x㯳C�i̻�eЃ�%�gC�>�@�BC	�y�	v�
:��CK9�&(�p�My��~_58��Vf9_��t��4�"q3� Ќ:�ku�]j ����["u���]Y� ���Ee�J��L-0����f�%̼��s1/w�}XYt�gA�ѶQr��G^�@�K��v���ɏ��W��o��n��3�?#̱DU���9⯕HA��]��/�čD�3{1�mX�{@�R�gF6nb`�� l�����h��F�1�|���2�h�^Dte���lV��]2Bh9��z�*��`"��76��J�������Bɔ���S�ggE��<o-�<\��e嚬y�����ٲ���{�	�|���w��[�8�1|���(ˌ���pT,���у���:�l,�],4L� ��A�-�SG����kщ~�D�%̰��gOWQ��N���ֽ����p�A�y+�ެU��Ow�:9�.��c��o$�j�Sj��D��
��>��ԩZ�'H(d�������vn��Ľ�q®]"�d�T+�"�[�����W	L�2-���Ďzo( P4"�AWw����_2	���EhD�뮶�fH��$nq.wo����q�g�W�zl�l��6=ך�����Տhѝ�T��qvʯI��$�(�2��O����Ip�J��15
�ל�h��d�+^-�نƙ+d؉,�(f��]X}[y�A���oK��"�z�/���G�Ɂ8��23Y�����%b���Ԋ��5Q{�c�s�J����>���jr���^���P�18�%~�1���xB��HR����a(�,u������y���bH�X�{O�{�����#�r��%��6��T۔���y2����q��y�O�9%����6����7�8�aY��dq��;>	�w9
���)�(�o/+'�����Z/�8k����1[��>6��Z�Q��[�`�2v�=T+�^�]>�{�ph��5�����!`��Ք�K���Jbf��}��&�׀S���&T2�*QU�tSl(c1c���V���o�3�c�S |mr�SD�Gc���`�tĝY�w�^�c�5a�Ƥų�:,6U�Z����8�������(�=���C�Y$@����G��I�䤂�x<��z��!���:	�)F��w�G�d`p��>�y�-`nf�@pWvj�=>�/��4�� ��;^���J���ʓ� *���uU;¦x�|��=��j�e��|�;��Fբ�jY�Ol_	5Vߢ�ŜXF��I��w@����Pv���=F�oߩ��4�i��(G������emG��G���I�׷"@��B��e��������y6`�A]~���^#Th�l�W0؉ʄ���Y�S��3=[��� ��]�
X3�_���>�j��#-l�lzz��&a���]�2���$sO�t�X����S�K>^���\�@�����m�SL�Xw�.%�UEUa*��^�GED�����	q��ZP���=�}:�Rήg��Y7�������J���18
�g��O`���ǤDG��`�ʼ��������ػ����l�~���i�+�f�S�Zp�ĺ���p������ .(��[�|�Ã�3�T�ۢ�#2�8Z4�5U�֘W�zڋ'I�`�\���+�wQ�$��8}��im��'���3<�Z��'ț�M�Qk���	�	�����j��7��&:	�Ggjb4�}]d�����"�����tX�(���k7���A��-�e���b�*V��,�z���h����3~�?��{(���e:v��U���&���ޜ�Sܪ�Eߓv��+u�b;�7�̦��h��QG&I����LQj�`�㑝J��[Fyd�w�A2um!��j˹rN���ݒ;��F9��ZTj]�ek&;��y��f�v�|k�+�X"���U���Ɨ	�Hp$9 �s�7r|g�0�����i�C���Ŧ�h�9:1k������p�F�s�}zp7Ʈ�G�o�H��|<T��E�e�O��%�{Q\t�'��es�D��VA}���L%���qsmU�	ǧ'��m���۩ŉ���W A&Y�CP2��J�'�R�O~/8�"�� �1�Zs �k��U��O3T�-��k�'�?]V=����_�1,�I���t]���L�pk]]�D.��E	���7hs{w�C���w��0�E��W{V��I��[V�U4Wm �	�Y��bE_��dU�J��	��KSk�cS���h�ˢE@Xߖ��~���I.k����c���#�La{� 
5H'D�M1`��=тN]6D~xcv4�&�8�Ҍ]r�/ܱ�v;�i��M͋�q�̶	�3�LU��Sʂ4z[�b��';���@����w:���gb/v�Z�n̤(��X�,�����Uv��#+�&ܓ�H�wr��-}vh�w���E*Z�@��I�j^n���TN�ms)AӲY.\��eW�O'��M�|�-�YK��"�<�x'=���-B����__f���th
ծ��e{6�i0��A�UfS;�Y�2j���m\�8Bޫa;������A&J��s�;��/$lw�b(��4�橲�.CG�3ѥ� d�kσ-�.�r�+ܽ���j��/d$����e�G1��a�	C���X���t���1����	s�Ϧ:FB+�\zOY�,��-P�o�w��#�y�u	v��x����N�.�&�X�x�.un��E��� \!l��x��{q^���𥸥�ޔ�t�]��[���-n�FLz�$}�SvQ���ďf�&ݛ��& ��R!��m-�V0w4��ķ����Z��5���OUߎ��f~/����-5��
�12|ט�#�9[W~Z0I���"ڄ��m�3˼/C�d���+$�y L���[B[JmY�P��_����=�Β�ֵ5�
!��u��|zܙYo�"�2aj�8^��hH�U~�k=�Ǌ�0:�Ѯ��f�j(D �7!'��Jw�St���ѻ����la�$߱l�ЀЬ��#�D`�lm�Ds-�րlyk�$$�D� z�v$�;_jn�FIL�oAi�͎���l:��q/x��\����%�M����v+���� fV|y_�|f��t׳N7M�W��?�Z_��?@{2����e��x��9>	Ҍ��"/�X���q~�&v�O+5R(P����mS��hj᭩|UU��dП���>���ΜC,h�I�xjb����>�3�Q�c͸�;�4q���8"�؋�xZ_��җ<ԯ���j�ƥC�?\�Q����o�p	(���I]�� y�gz#�^��Z�z�Cd����-�͘!�M��7O�ά�XI'��%�QqC��A��fS�ע�����VbL]�m#�.n�VHȞW �:>1��_�Y׈���a�2�_�u�s�񔍹�������>9T���}ep�KHzZ��!�4-rTU"d����>8�s����,&<���gQ�����-�q�:9s�`�`sV��?jM� �JE��x�p!��(,�w"��XtRx��T`���R�$�a�V ܳ����ڹ]�`U�I���VX},���{�D� �Չ���h�=�H��R�vp�Ʉ�'vf������#�>�����}��έx"�7��/?�"[Q��[Z���2��Γ�U�a&��(oA$�qхgZ岜�B����<s_:�68\�y������~3�i�+�W�R�ob�F���cY��GS��������P'�c���L0�H{��{�YC���$����t��):`a�Rwn2>�L޻/^�]���,����)����N(1�j���{V0k����/�\N8�@}��s�B����EQ�����أ|�M��%W�}ȳ�Y'4~ΰt�n�,�8���*[{(��	:BT�߆�u��+̀W��s(=
#�V*Q8��+�Ɛ�k��E����j����n���Y��G�4��y0�����'���I��ø��I�q���MTS��+�;���\DˊE��ʕ��'��KNHa�� �7	���J$��?c��ɒH�ق�A*pD���^k/�^);.�Ⅾ�h�A����9�N�S�}9bҴ\��� �,=��]��ߊ���k�=��(��n�ю�sL|���R#'�Pz'3+��m4He�6���)�-:2��/#`sPs�$T�ֳۛ\;d�����¤ɀ[�"$)BR"�vO{,���;�n���v`����"����;Ţ��r	.D">�'�΢l!��c";��>M�S�-K>dW��