XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m���iz�A�Nn�h6��ڶ����
�~���؊���%���5�|�i�L�iflo��	9����v�y�V"�ޟ
U�4n	��Dp6��\��o���t�h��#c�����ϭ�<܂�!vHANY[6���xm���K|��pu�F;8�ϑtG�Σt��|M���P6�8H�сh��_�8a�u@Vh853?���>xd���MAw��Ay�,������y��%�˫Ж��bR��� ��*z6eٕ�1KɊ���x�]R|�CWI)pX��2X��Z�w�3y)�\4;��,h��y��J����
�;(1�(�Bn�tvr�J_gKQ#��~�!�=�]�{����px��\-p����,���L���Zo"�׌��DZ���ky+���9�]|:�K�eW7�� b���������L<"`0KN��7�)9�H���\�.n��g5P�9(S-V�3�:}��lGpg�8��ͱ��Ѭ�Ŧ&f�F��|��5��Zã��M��󥒅��⬸"
�H ��
E-�	8Ju|���bƲ`ș�Mh����e�����kY���"K�,� N?�HRc�{q�������_Ҡ�(Z7�1�p��"� k��PC��|V�U6a}`)�PFsUV������"IP3o���*m�J��]��s�%Gֹ��u��𤐦u��٨�!b��=U�_l'��՟���D���)O��������%�FJq�d2�CNƯJ=���X�m'3֨�ǜ:A$��s+��XlxVHYEB    1b12     8b0G�j�������s�D�O��>:B�d��_��p����Gca�9�=�1����i,�Dk0�h8:��uҔ���=
��h��n@8�k)�g��g@�����c�Jˋ�$�z�����ʌ�e���<�`ⓟ�9�7�pjv0I���3����}9�ɲC� ���(d��MX�8�p� ����5*�`K��_1<3x`M�?�	��f�|����p&΍��=}9����鄯H/�q�k�T�ya>���ee�g\�`z+r��eJ��@ӿ]U@��aS<�/��%|�����+��GC�݃��Ke�A! ����V�a�Ŀ% ������*bs4�Ti���L��q�4l�o��;a'�V�N<@�&z��5l��+���#<Ź�1v.<�8f��]?��~1'�h/�C,�A�40��aw���kr�x�I�r������o��}+l&�s!xD+��9A������������O�n�OyB�d�;X:��{�M=Y�(r�#>
�e���=F�)��ƻ±����w��+��GJ����	���_7=���}�N�� ���׈f�.�^^����E�#F�k�\p��B�r1c����pQU˜�
9V!�F��SgR��޿AԤ�R_"���s�d6���mG]-��<EV��dA�bF��E�����%���3#�uV'��(ѱ��)g��1��Z#`��M����I"�Y��u��aB=�U}�ɗ�؜?_��M<p���sH�#�ARo(
�R�����	�\����|E����p���-l�$�$<S��r��O�ަ�9�8��SS�nc4�
iw(� ����#���g�f=-41n\sx�{4���C����ҍ��.ӢP�Ĕ�DF��[���qYCP.�L�)ݏ5n[͑���浦>�R�����ʰh<��S��7�U7#���.0�����a��������PGt����MXYD�KVM�N[ ������8����6D�R]ֿ*��o��"�d���6^��{741I.�݌����"Dq���=ĉ��X�,(�tb����(Þ5�����?(ѝ�{�6���1�E{��7�j�����ȩ�K�s�.t���YO1�faS>�\����S����,�F�)G�6������M�/�B��/kSu���	˝�'�r�P�A�s6��4�;DcKi'Lu�]d�3�l���y�_2na�[)��?PV�m���i���8���e=AM7뤫�|�s"pQJ_F	o�b�9mUH��_��V��*Mb���8�aM��*d���P���S�"��\���IL�H�K��[�a#P��sK���!����4A�k�\�N�\��Ҁ�W,��L���S���Q�nF�}�11P��4 T'�dE���KL\�E����ۡr�֒�TV ��I��)nǦ��z�K3ؖ���/�~Ɇq=�?@�����x�
؏_n���l�R�;�M`��+�B���(X.��3��R�d^����-���i�s�w�?K�� ޽�{���JtU������� %�r��I�V&\Dߝ����2\�W�𛕙C6��~X��=A&g�qge����|�Ec?��X}Y���i�"�E!<�X��
ޭ&?EޚƖNHeδ�V>\9�
ѤY��ͼ5��\p��8n�o�6�d%��6P˕$�v�ƅё̳%��㎳ې˰�� ,�Ҿ���ɤt�,��b�v�
�`�Ԙ���	���r_Ov��ae	�ގE=��Sr�XR�5"�-���KP����IF�v�ۆ�hSl��H!M���F;p(R�����-�ch�# M9P ����s/�"yw��oa�h��$�l�}�b7S��H_��d�ÿ]�HH{Ds;�ց��p���kE�\��������ͤ���D0h��|��� ���?h����s��r��.��0�,]���+*��uR�W���Q)�}�kԝ�J4Fn-ɦ��V� \�l����A^��;��w*|Ll�τ�r�'�o=՗��0�dj���%}�����0�y�ǔ5$O+'�h�����ۗ��Ɠ�}��SBw��]x#�HV,���r<��"ԡ���$;�X9b�ݛ��U�TB� ��������A;as���!�cjl�Q�c�EP�t�G���{o�4.b��F��"��\�Y��