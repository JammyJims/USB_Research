XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p�|��0�7�%"��!�??�]CckW9*���+b6`Ɍ������]Ur�1�Vs���אqT� �r�U|��D~�.�s�[��YiP�&�鳲�WVe�(!��m�~]A=��q!G���ņj��De�*q0;9M��Id��z��x��%4N�~���-:�2Z�'9I��z����2y��a�93+��Rȱ�,�x�H���}�ԓٜ�;�?de��Sǣ��xu�<l�o nG"e�����.%4���Rr��
�S��u$O�*[&�@��\�:���jn(����OU��y8��e�7�\Z���|�	.ׁ�mn'Q�v�r7�e�	k�@T���Q6�X��N�k�ؙߴ�=Sp���y�����Z*y�M6ُ&�TW5*�٭%������]�Nz`�	NG������V���K�f_��	��#R��p��웦�`�E�9�>��4Ii�V�h�r�L�?3�Kτ�\|́�5m���X�zw,1�Y����@Q�ۇ���x����r�ж�c/�2v�")`˪j#c�'��½Y@�`%�E��(-ɁV	wJ&���Os�r>��J��Y��K:>�J�ox�BB��
#nzu5�s��8*�o��7�MD��3�@h O-rH-�Dm��Rվ�������2.S��HT�� ��'���WQ�����@{qZy=K���
x�2]9�&p�Re�<%�{1�eS ��U��fIkݿp����\d���2�	���଱v�$,M��P���XlxVHYEB    cca4    30f0�kF��f���1N(�� '5�;N��d��p�Eh��O�?�n�Փ�C�U/�L^�g.��ڏ�ӵ�����#U�b�G��^��X(DSQHP��h�ʐ��l,ߒ_s��4,�)�F}F�꬧��U����۪�1m������ h��j���j )֮ �tr��{�pI�E���A��A�EҨ��H\f���K���xG&���}�a\�SX���8<�c� �+���0p��J�h�^X׃��>4���*���s�{[�PA��5v�g!�#|i�\���x�r$�L�%�aN��L����%�Ȟ���4U^��(�jd���d:N�`V��O��i���@d�x�sDk��c�GXl��l4�~�6W�%���9��\��?/��d���,�ɯ�y{�\�������Q��8�ː1�Mt!��}�D��\"���v������n:�2���q�H�o�kyM����q,M�!9���? ��"�a�b�&��(~�K4[5bـ@�N޶���Zq�)��mR�n��,����h�=a�۶�fq�k��V�?P:�9�L0�7ߑ������ا4�#8%�⊞¡����ӵ^�����C�=L����LF �]�$0��eV��9Gak�g�PRr�[/���Rh,%��L}P��n�Aw��X{�H����X�4d>���L�a�~>��wCQ&���^�%T�� ��M_�C�%A���f�Ӂb�ڄ9�џ����_��F�����4�V�F��#o�Y]Wњ�F�f�"���Wu�A���=-��F2��eh���1|v�:c �8�:�������#1�����jG )7�;��i���	�*�.��y��c�!ɴ�%���EnU`v�ħ*ɄҌn�\vrS��#.}_���]O��d��}#�.�'�9y
Bm~)��a���(�(2��7�����ly"T�{�Uhi����k���0�P7m�O4K/�R�wd����ć���{����tjdn�_
('m{+��dg����Y����i�N�S����&Ի�/t�)8�87@�3�|v�!���N	�����KG�'��o�x=�Mf�߫����̧4a*�g��{b���r"]���A��(��5��m�H��@	��� ���~�]`??�fz3`6���Vep[6��@���|{t8��q�]�V�lڵ�6���H��Y򇨂�W޻��
+3�.��TY�w�T�����Y
-n�h��b�R%+1
�ejI1sܳ��������0W��z��� O�a����O�����aC��7dK�R��x�EJ���?�������	���Ǆ�o�V q������ڿ�M_��s�mSS-���yjP�ǯu����'VSn/1�$�ɯ�N�}�KƚI���>�eNC2��
:C��KG_/;�-YWC�j�&�6���\*J>�2M�*2>�}t��D����q�e��G��Po�K�!��FTY�ϵ�����oS-`� ���ɩM� N�m����=��P��|z@4.��{SZ��ᷟ���**���Tp�ѓ�J�}��@	�R���D)�N<�����Y���}���S�m�`��UZ�v
�A�'w��ډµ{��O���,����];,Ձ� �3aU��K��:�
�!�1�q{����\���m��������V'���I�y-\u�4���Q�4�f��k�0�L�	ӚK�_jM�
��j�Kr�"��,�b�#��9�jz�X��"�K�Ws2z�X��'ŴTR��e�<y��ձZP
��'�)�H'N���'ՠ
%���i!��mRq����WVr/�t�dJ�Acn�g�C������\����s���c��g�y��`���"fq��������Y٩���!�)R�s��o�ӴJ�y7����|��K�\B�H���xT���o��G�m�5]�r.��6[����S�:��t���?�,?x���9;���|����(�F���c!�d�7�$Q�����p�d?6�솆*M��c���a
VN�����cWeڎ8�p�F�V�.�7r�7�;�_62���*=HK�L�+tX���iV8L�W/AE,m�$r��"Zzj���K�{��,�B��aLO�:`3��I`���^:�u��:���s¾��$���g�. �b�Lc{��}�W�^%��Muq���fxm��t�{(� b�W�8 �\_���/����ߪc�q%�P9��D$J��}fp*��Q�d��Е�`b�ia3�C�0��9O��	��W^���f����vjt"0+,-�!��y��Z=S��)�� �JbO \v��Դg:�+:��r�z�%t%Z�YF:^=Y|jL��@�t�D�e�B�������#����Ca؁�!�C�y;�@�s�M&�:��V�	�Y���{� �����c�{��כ�ݳ��1#exil����3�{���^!�i��qy��i�}����;�������|��&K��U�>ܟ���_"^�x�d����C�<2Ћ�Q�w��k�dc���ά/�4�)�P?tSȈ `��r�t�tи;�:����bm���wCVH�#���$��smp�A(����7�!rr�~Kp�t�ǂE�T��M��m�(!RrYD0l����%�ʪ$P!�)�ך8P�PL��4q�����1����7�񂖱Z�R�k^�!3$�b:9m�)\ڵ6g�<e�d�Z0)~�v>�պ���T�`ය�㏂3�7G�����Qe_H$�:���o��A�)?�F�t��6t�7+�Yj�X8r��ܛt��:�VΈ�cB1��u��ηܵ��,�%��]�����-�f �Xy~���]��)u�
I��Ό�H�����uL��>����`�*�& �׭�vCo�T_�2����@�y\:�)��.�ة_���ꭷ��v�(2�%c�y�ƣ'���w�R�1Nw/�6lP>���mEqy�������	ZR�8�-7|A��,>3p�1pnZ�o���(�|�XP��~m�~؍��F�I-����dҾ�X�l|�	R��K���ء��[��
�r�V���@���'�HYH��en9�-Q��X����lvE���J��떓�S��J���� ��t��P�Bo[Ƶ�� +��*�a>����-&��܉_|�D��D4J����&]�L�[E������l�X𠱩ۋW�RSU�e�tx���
�4#Z
��h\yI�s�ܩ���OOX�b�@b�Am�L�R'��( ��8zช�2Z�|�yMS#5B��9�*e8�Z�}@{坸6���&�5c�!�����s�
�`�E�Q���E�jly����i�s�h�ʶJ����+�QÚJ��;3;u�hyY��O��Dg���
�{��j�F�(U��B%�-%����X��"u:BJ�D�(˥V��fD�b
�!	R��8����Om4.�8Z�-W;�0R�I�g������{?_4?5�����=�B�W����v1��`ʧ~��bIyr�,f��q�M���\ F��VhJ)�zPȑ��9��I��<�D&5��:`J
���p�]��" \~O�܁n��arjJى՛I�f���T%��gjzC��5�JYϑh^���u�ٵ�s^�*O��^���}^���us�n'a��io��eQ`�$	�{�.z q�ݭc��#�j�?�t�/�/C �������"{���#T!�:�耤�_b�w�L��`9��:7�8~Ƥx���C<���i�������H��B�s��q���q5^���5*�'0�*5�'�a��y�4Q㭎�����oX��UaMR��c4���AA3���p��0c6��HB��ċ�.�npF�&=�/R��.���M�;�T�Tq$nL����?�3�k�>w&�04kPD����Z(*�"�F[�V��"��L�A��A������վ�{���RHN�nD���⭌�տ<G��W���愮8����1�H���)r��9Ab���8�vza����\����y�[0<�8R��p�
�BK�A�ve'��d:F����a���8�]5`?f;j�@�6��l�]]�K�sl�[�.=t���/�=�E]�!7D��y1�5�-QI��X�]�Q��{���	?���X��oD�U��R���m��G"�V\�{��!~�d��6n+�Xy|i��J��8s��u���V��C;L|B^ޡ�p��D<��K���h�6��A�InP!��u5�C�N��f��+�E�A�w��:Nk7�S��ǰ{�&���}PX�4eV��W�:����p	B,�/���V_���}���F|`���Mϖf��iMй�ұ�7�jJ�+������3E:H[�Q�H��!q��Y����P��x!7緶��Ǽ����ɴ���6��/��0���ʞY�//��Y��ug&hUD���	6=�!:8�K�[�t�#0GPq��JA>xj���)�[���a�)FC�љJ��v�m���'�x
sC��X.
�>a���C��۱�������[X� �*^*��4ϼ��bz`�M%6�!μن�<6�,W�q.:�k!���ƈ`��p��8�������S9�H�ʎ%:��-/v\�(8���gG��AP���P1��(�D,!�w*1A0�s�;��;���~����2��D���.0ܹ�(qL��]�:g����\)���#RLw���]5��Pg)�I� ����R���#��_�t˺��[��(���Z�,��9�ϳ�&a���`�S��6z ��|c�̮hՖS���G�Ns�b�/:��$6���\��d�Q��e4��钁�n:�m�4��N4�^7��o���:��Lo�}�g���y�z����̪�%������v�d���N� ��*?��'U'^�֨�ie�h.���S��}�n�ݲ{��%�#��-�A����"HWfH�vFL��� �@�� ��'9o���ߌ�=<�'��G�B��ߤ��tYŝ6M���:Ӻa�\���� G��(��= ��M����CoJe�AS�v�� SSG��VeH���Tw����6���V�Y��w���_$3�#J�MIb�l�� �NDg�}	;�>?�KK��zG��%Ǔ�Z���锗���_DX�Y$���U�s�ЪS��t�hl��B�'(s
O6� B�`�3�Q�j��Q3�,Y.Z��{�M`ܷJ�!2�x�3d�z�'���3��I�h��i̅�'V3�����pA�b�P��5�q�"��4�|�f�dr��?��iʠb��N`���4w/�G$I`������L���.�Y��P�3�Ep[��[��bJ�+��v�X6���̮��Q���_}��O-QNHŪ�<��;���k�E�q-�q�<IW|�~�n���M�WR2t$O!=a_A|q]�G�+��C�w)$��6+� "��q���
bL���Gl�Q�$���B��l>��u�e�\J��}��E򶆸� [����Fy�UX�I��m%����B�LE����9;���~�����s3�ZLuXj����Z�!�rI�?k ����$R�yB�F�=1Åӽ��aŹ)��@��-҂��*,����s&X<]��e�.�s�G
���fǒ9~�%
��=:���8��~qaC֑/��>u�1:��=�|j�s�Gn-XP��A�zA�D��I�{ P`�~eG�A3�X����h�ɛ����(�%������bVI���"��h�O+*[&���#jO8�9+9-%~�ݵK��*���d�%g*0�O�dc������ � ���^g�W6|$�d {��xA_W���9������:�'��ũy��������{QT� s͏�f�t���v����F�q��$a%��f<�j�&V�.M��Gz��K�Z�m	&ܜ���65o?�)7�>dO��I����h=�U���v�g�l����Ŕ��φ%�qa��a�9\9��w� F��w�j��ć�A2��dGuw|>J�Mu�&Z��uƜ��n$�N��̷��w:�6�����c�nq���vF����/�詚�?���󀔜�����(S֐"�2Ҥ�N�����J���.մ�)ۿg����1�5eC(�+kփ`����%��.�	��{�Ů�/�W�NF���wʋ�D��~�e5��=!�v�NO�܃}�� H6>z��?��S|�y��A�	Q�� 5���u>	x��ν�e�<U�6ɡ=�eH��صz�q&��$-�����Z��z?����%Í4�ڌ2x�����-�``�9��/�Ky��k$�v�RJ9�������ui�3;mi&��t��؎;�+�f/�+k������s��֔bP)[�E�E���G�a���>���������A��f�;�u�?����L�A8������Kʗ��5�y�0��s�ԋ��(FS�s�; ��]���
�wr7���~O[xf���G�y��!��~��Pnc�(��?����a�(�T�E畩W�4��s�b"(y�,\j��^������佃���'�y)���$yL��P[��5������FrɅ̮��"�hͲ�'�:����u9��K�q��� �sx�cHD�<!��P~�|��P~S6(®�ym��1֣�
�R�v��lPF/x��n�������V�Rh���˦v�j�����(�>�4M�o�w�LJl���a(+r�� )�>��@Zj'Nu�`6�\hT"��quh]���^
����-��?����:��MD�w��6Q���M���
1�zM�7Y}N�t��!q8�pE����HQ�g ����6�(g�w��v��2�׺�GA�º�<���џbQf��sp���P�%K�x��'�D/�q��`��wY�`@��YR%I���@[8S�ׯ>|C4���Ti�:��������S#F ���|�D7x��TՒ��X�:�d$��x����}�.�3]C���hT~�;1}�"^�\�8_�w����ɨM�������M��?4�,�>��hO�%R�+��1vc�������9~)�g��È.����3�P���F�o&56�&������荽���J\�:ɔ��cǥ��8�/v���q��*�ӑș=���`N�'H��0{��3pOH��ߥ�)�H���Q��0��|�	�vg��!�k��o�`S!u0RT�`�u]���}�4�\p����CjH�rnp^ݽ�
���ģ\�� ��EəE1���Au����m{+�:<����4T$x�~����<8d�ۤc!�����J|�l���\�j�*��[�E���?.f,�Fl��?�2���	B!���ŠB�w�S��7Z`�w�Kh�,�K�*qJ��S��RպN�$-o3����e�xw���۲�O���IG~����a�WK�9t�b@�w�L���TH5�"�}�/�IM!]�*�G3-��X��e�Jӓ��b�8� �͂�q��z�]L�ߥNM��F��Y	 5�Ю�j�Ȱ��f���]���󝭚3 ���z�4X6.�I~[W&�U��҄��гm��L�M>	��^E]�m4�'v�����BK���8�����Uys��j�ct�\#�͂>QǍ�_t�MWP��Y6���oh��P������3�Y�uy��ޔ,Z˳�M����
�h
�|���U��c��z���#+��ґ��/�d9>{2�B�F��'��4��3��Yd�TU{�)jx��<���s�AU�MJ�,�4b�0Us��#{��@�v݌y@C�$Q��=��5�W��x�4 �Y�o�nfb�ι�?��T�z��|���a{4��.��%��R�6V�Q2�Y�/���gQ��=����r� 7-��Ӳ�y�f{���(*�Dt�Q��mvI����=����}e�OZ���'�Z�2Uǂ���i.eS�}�/�Н<�"c7_B8Tϟ%���Bo��\Iם�Z��p9M?�rf��5��z�5�=��0@!r��W��?Cq��Ub�'���pK�?+�r�����ə��x�5g��df��B��e�:c>�� ���/�t��ws���kN�P�\�h@��UCX�T9a;�q_�v.;33����*�n�V�A ����Ί6���< ���K�P_s�6��k^�\�Mz���[1~ !�7��`N˘���(^��y+��y(E�!�<��`��;�ʲ��������Pl^D��\܋ů�,����R<T�=��?VK
�{���s�~�r�b*6�٩>�j�.d�ܠg���H���g�3���ņ���qD?�KY��G�h�O`�T����ur@2���%��X�T(p<)	P]�ע��{2~�0�G�0v@�ބ�1Y�N9!*DbBq��#�<ۣ�fE)l'�(��tl���|�q0w���*B�63'�DM|�t������1���
o���;q�����E�M�.w�h�h���7�k����=���L4��I��?��f�a�	"���2Y �46ߜ!/`��Hdq�4�{O����W�e@K�S��a��-r���&�]��Q���pxc�d�����ۑ����������S��F5w0�,K|�)1��-��?��YV��IP]1���07�,P1����?�#�9f7����&�{���D�yq��!�r�68ƵYt&��y#�����@����;�_�| �yɒ9�h^�2�޳�
qt>�$6|e^ء�+������<���N7���K�[����2�n�������Y	�i"��\��Ea��M���*�߶��O�詵�I�D0����w�v��Q �y(�s2gP:���^A��ȟd$4�s���[(BcZ뎪�X�kK�$}���"�c��F���G�*����H�M�y.����Pܔb�7�F��-�F�;�o������BС�*�
���7|������B&�~P�f���p��p���^�|E�c/*�:�o�q�� ���r�v�CW�Y�k���u��[���U2�%��X%�E'��߰^�Wrq�Ay�Q����A�������,�,n�l�S��^��Rl��o����'����$ʟ1^L��C0"t���Cx���RMNj9ϔ�v�8j����X1�_hD-l:l'���p|���ca5���B��*��ӨK���r���I�d��
cI0�=�_�t4;>>e�J��*:�[��dL�[��A���D�/��<QyE#�ĥ�RW�c	H{�u�R\�8rv�S�'|�B]/y[Ta�ż� ���:ۆ�ڷq#9.5��$��C����d��C�:��k��)ja{��"� ������-����N�or��ȝ��. �W���_�M8a�S���W�]O����n�~�ok�?2v�Or��ex|X��&`մ����/"W	Ӏ�O7d3P4۪Y��$D����P�؈<����"���夷P���S���&��,��u�~��\{Gl�~[��-Ҕ5deD0 ����֦p]m���^�Ju���Is������8^$At���\�B����>���e3J��3q���q*�Y���=Q����e+32dȃ;w�4�7������FH�@�J,�wr�����:@���� }Û����	�WV7��������a��q�>�f���V �8�B���f�) ��8��<�h�Q"*������{=�k������.DY������_L�gW#E�Yi�#"�I��U:)J�b>�CT-�JW;ɛ��凍�%���Z! ��8LjL��J��S��v��&X����Z�E#�/�d�M����=��v%��O�]��[���Y,�;fA(�E|����v�TLtWO�7bׄ�@�6�c�4Ê09�?���O(�(�	G՗"�s�Q�����N#�T���p��D���]��h������|�ܐ�_3H����GEj�����J5���Ӌ�3-�� �5�U�h!���wVaWUuժ��W@�����T��Ez(p��&x�L:gn���)��'+�+@RFH�p:�#.23`�N����7�WѸi�B�dckE��L=�xQ�t��MbX#U,2�Ą�|\P�M�"�n�����/ip	g�g��@и��,u�pcl�g�s�D�{C�o9�JWѳc;2m�UՕ�/)���2�\E�-I �wC��Q��;b��(#l�w����6
��L}�&>I�3�E�~*f�������a�{�v���ӄ�]]�Fv�Pm��l�9;��ZNr� �b��īܟ��N�Xu`m��^�(���)u{v����@	��.D���������Y3�h�e�Jj���{�!R �8�x@�$�5�v�T�[�]���#L����功S�#��F�����4���h޿��8Z����|F����F�7;,pvi�گ��j��"?+S����:�q\X�s�� �_S��2���ӵ�f�ه�!��ԏ#��#;ˈ��-*L��Ɏ�'�����2:kP�cLP�ô�T��oQ��G.�I�9L�nϾ]&RQG�]�0�F�Q٪ex�	-+�y���աh�|G�*�Y����cr�*���($� ��Dآ����x�O����$1�I��XP}��M[��P{:]a�q70�e��ՠ��L�����כ��d��T�Y�������(�ƨ#�/�wL��c6��S�7G�n0����-��R�ec���5Op�V�~w�X��Z:�m>Zӭ�0��4Q��_T�J z���fm_�I�W	����8N	�G��O4{��2�( R�������M��&3��ADqMg��`G?�\*K]ȿ��v'l�WT��z��n�C�ν1?�]��{47&5Ÿ�X��Z�� �1�h��G�e�����ӄ���� ��1F6:��5�2*�������/����ȕ�8S)�=+b�Q�i��p��8h�r߻�Z�I����E(�6�'���3F��)�~=�7������c=2���""Q�����̇���Ἰd�������l�0&�p�0$�e��¬�w�{� ������lI��j�m҇�l^��[�#��\�#���В���QZ�=}ce���W�P��5�$FvI��w�Ϭ|M���%�O��G���Y�lp�qr&n�k�� ����c����l���Ύ;J(e$�|)�p@TP��fǱS�4�#����U �s&Ĭ���ޒ��g�	���GOY�4�A��]2 ��=]���.-*f�s$۫.�{ʸJ��d��?;6���p�y!����Æ�:{�q$�e�j�d-��8y�ЩV�7�'�FԲ�d~��%|ūg�G��Jel���ӱ�N�lXi8���]�aD߶��ۼn=O�Pr��at�[~�+w��'G����J�z�fּ;E��m�}����#!���m��w��w�	�4#�*A��X�ص��։gC"�ᗂ㛭����/9¨�;�7�
j�n�o˻0��`�o�Z"��
�U��(�溆�b��0��/����5a�^h���+�>H���)��֏���,l�&M��e4n��P͏��vL}���!���c'�-��Y��+	6�H	�Y;���L�z �&�Ă�`�8FT�\c������nmƧ��^�7-O�-f�w�I��V�etj^0��A��x��ՔOR��&�ʫB�+^�Z�D��f~$װ��Vlk!�����7*�NPW��pK����?ZF��H&Htf�'�B�V1�`%�Gt>я��Meõ1(E�HM�����f8�VI��������qX4l�Qm��h�3��j>kK�O,�3��w:Ԇ�\�֬&�l�f�se�[ �Aױ�v���kz {~?*�Χ5�_�w[v�{ ��Pѝ�m^�<*�L���&��lx=�F�ڷz��Q��Q�
}W�MGzz.T�qS��t�=>M���2�X�4��LR��lkPݩ�.z5B(��j��Tֈ�ŝ^��3���]"=_����	r��T(�g^`��#}��kr�+���.y�=Wюw.��lO�$�cu�,�/q�.�;Թ3���"�E����8�ǒ�����5	�:�2�X�|���X�v��64��ՅT�Ot�[#aq��8�^���}�5��j��.��XCC��wR-��a`C��`p�`X��J+�wP#W)1�X($`!�N�~}?F�pfoX��*�7�NXՂN�Di�\���7�V�Ζ�g�|�e&v��a/*c�(����}=o.t���zg���ͫ����h�F#�^�P��c`���
/_X����&��Ѝ>� XϖR�5C./ �%�p*_=G�vYpB����Eo��|��ND}���7x��A�)4�M�'���4[��