XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4`� ����dVb^)��h���rߊ%&��8GC]�ђ�=�T'���?���?=��D�t���5

Ր�I��?�Y��qS��%�	K�K�*����.�l����#j�l�%0B�Q�4����n�^:��Yvy�5��\2}��9��n�1������.ૂ�<_�Z�B�K����sqnc����U���0R4��a�z\���Ѓ��`'�<m���"�Bu�����G,E'�R��91�*�������C�3�U��Ş���µ_kz*����ǻO誦����T������Z
m{�ѱqN�û�ѵ�U�hQ��=�3�p����.[�V1zL>O��qS=�G����juU�Λ㻥���F�w��(̭Qђ�#��7��\�q�G@W�B��	���FP��JB'�6���������;�(	YR8"�U��z�X	8�[�2� 9�={6���|(��q�c��@�?���#�>.��e�S���x�����)zd�w���dR��W~��*��z��n�����T��_d|�OtښӠ=�k`��������!�m�Af�w1F�sw�em����!�B4a��8�V mk��#������;�Jvl��צ�o���C�ԗaY����_ǲ|Fd޳�&��<#�a_O��Rق�UB��z��>h ĺ��OC(c,����{��Ng�~�B_���D���>3{�ߺ(�~����'�tɩ�w��d�Y6���ݳ����š�iWmV��%���]�����xXlxVHYEB    ce24    2d60�I"����jX�\}�55k�v�-��R��$�a|�
Z�=�/7��7f�r�mf^BU��,��UE,��;�E���"��z�
:�6{U��YhF��NR\VS*�@ԓ7�[, o��:��$=�1����&Hx=}>om��j}^�șt!v;y\$!� �)�� "��꣝:�itR �`e�MO+��a��S�aȰ�!<�U֥mO5�
��
+Pr��ܜ�� ��Z��ACq�D��y�lz�\F��c�N�ؔ��S����Zm(@޶��pw��C`�P�rR}'	�ځ��x��ش%L8�j �MN2���i��0$��P��4��*�5�+�_M����	���#HU�'�U�}��I���Fa�đL=�u/�h�ap1m�8��*z
tXl%�x���kgagM����m�9�V�H�����`�Ql#����\UQZ��Ȗ�v�ڜ���Y�>oRޥ�hlӠ�e��}l�W$�pX�Ǳ���F
�qa�q���$x����-q�b��V?�����X蛆-�4p���G�k>�q�d����Yݮk'UT��)n��J�J�?X_�M}i&��;)�z�Ww���'�s5��8\a�ؠx�������g�6j���9^߰�Z������Ƚ'd�u2/��c�-dv�uč��݉PJ�,g�"�rs8J�vfZϡ ���t[{/��1vxf��:Bx�H}�Y��8��Fn(%|!󶨬 �h�?:/&_)QS�a�n�A-��e�0Z���ɼ͋o����� 5�ɺ���r��8�>t+�K1zo�J��A��1�X�Cx� .�P�:�{��<����� w���4Vv�Ub�2��+��̂���t�{��rYG����ٶc]2����0#�d�.�`l{�*�u��}wl��(��k'á�~7l�[�	���-�?�-Ԃ��<3}*��Tgޯ�r��<t"-.��բ�ˇ�6h��Y$Y>V���f�}���9j����%
Ӌ�j��F;�dD�8 @�D��~�q��V�P�_w <��B(�����滳�+ s,�<Kx�l~3��x�I �����@;�3����a�e���t����&^sD�u��
߃ղ�UY���w�,�G���g������#��Q=+�W>V�M���mc��'�KrWv�[=�~j���W���;�D�ԊY���5F��Od���LD'�u��r��(GQ#8W��e���<f�,�*�(m��l�������sK����u�Ö���������8`L��WJm�F˝C�Ȕb�{-���"�@ ��j���L���$Qzk�[�i6��ԛ���~8ڃ2��t�~����,���֚�0���Er�.u*A�I�Z�>�k�t+���	�N$��S���S�t�9��]� ����[�q�[�U�^/��W�Ҋ�W��e�z��T�f��aΝ�cF1�B�`U��ۃ��KҌJ�zAy��B�Hth���4§�}U6�7�L��;3e�p����nT�V����#\VdX�.��A�b�H�Yj�:��3��J!��O�n���l�%!����q��v�-~����/f4���I�� ��
���}C�X���ð�ݩ?��xrw0 ��v��̄XyrԵj9���wʵ�яd�뽒.�@4���dq���.l*h�b3�J@������u�g��`�h�*1_���q������m�������t���Y�����(��P���bSM�h��+g�ʱh���÷Ԫi���AΦ��tǶ�ip���u�ͻĆ�Y�i�s��>��v�Ƿa�h�"3�"r50�`.���yW�)��YG����Q ~�Es�<~���h��d�M7kOk�ew�[���f�	5�u�GE��w�Z���U�p��Raz~��,�|s1��w��.[v7;���I�4@iX���Oo�2A�<�2&����sJ��}�V�O�37��"[9r��Y_��G��{B2�|����Q��S�����DG�V{T:ʰ	-&1
UI�|W۶c�����6�#��0��O�������r�X;��l$��Ӂ �+$5��v|ԃ�ۀ�u*z�L~���F��gN���6!�-���N�`�3��)����Ϩ ���ס�&�4l5��-3ܞw`�/%�+��U���߇މ�ǧ���(R��w��r���jĝ��qq��g��^>@����P�
�*D�̂������!��Eً�O9�MAJ�=�̶�'���b��O�	nQ�8i^`�w�˶��G��R%����b�U,SL�[�+^�
^��N�Y�)3�'^?��F��;ؙQ�~'0�?9�mSH�"T��M�ۓ�ª.������ �(�C�1��Ю�8����"�qŖZ�D�����8*WCw��c����h+M��M���+��0hC���u����p�a���4vE�w}��?�	���3�^j,�b;fS{���*V-��8��a����.�(J�,밅��m�SgN_��e[�q6��d,/"���*�H�_��J��oU�����r/'���6�5J��%i>�6L/�g禢�C\��̊�;&i��gQ��%��/���7��W?2����Ԇ!f��rF :��x1��Z�PC��2�O�XGT��lG�v��_|�0�/g,��t���|ا��\�S]��6JWF��?c:�~����UXDEz���h{�������:�����]A��zt�r0����y���b��s��@��aP�uv��!��(]#�ց�+���&'Uw8�*H m�^K�@��.m��xMZ�Tj�%QXS���93�,�9{�V����-�l~�Ǵd�QHڦ��ҟE[�じ��W)b�Q��$�+���F�R�.F�o�w�ֆ�k��Wm�_H��&����5ZR��-�K��~�UM�F@�����v�J�I�x�}k�#�q�a3���Ŵ
�"R��DW��7�b}z��Y�"�1V�D�H5������IR�Y�?~�����hs����,)8D���nB�@^��0mr��n�d�G�>�%OU��e�ڝt�d|�t��׆�'�7w�	_�Ģ%���<gkm��s�A��)q��$��k���8�a��h?۳�����b�u���v��D�E�.�&9X��Ay`f���y���垌� 1)�c'��?5nM̧��'d5�G�m*в	r�$i�wh���!�`ߖ�o�(L�!����l6r�^B��h���q�����%q���� �����$���~p�{��Ep���Z����*�9���K�j��lu��Ug������)�kp���B���H6��\��z>vs�Zq�)r#]�����FB ��tM�%0/S,��d�6k�ۗ�|� �y�T��U+��BЖz�m�S\��
��/�m���� N 섶�f����<��f2������ݸ�%�6R��Z?ׄ{�V�\�>�vڥ����yS�\D�~��\�U�X�״�ʍ���#�XS�xS�*v�8�UI�'a�ZU�e� V��a� ����h�EL��p!����(���ݦP���5:�Y@�ƚ�z������!Kn=��i����Z4�\E�^��\|�K���8���5/��]�u~�GJ�e1�p����+>4&���eh��ӯ&{�� v���`m�SP���mr�A��q������x8�$J#x;2�t��ɲ�Ƽ��%��]�=�=�zU�h��E�������#m����@C�%��4�v@˂�`�O�A5��L-Y�G��J�:ñ�|�qYo����	f��,,�Ęm��H͹�����.���:]����{�i���[���˔��~`�}�<K��Ξ}�'�!��B�zZj�%��{��(�*\Geɉp�|���'���#��N��x�O$�=#��^cW�^-�xL�ʹ9-�S-��*�\�YLA��̟63Q��Ϩ`��t.�6��q��[��4ת^cE߻��X��hI_�.1[�������R�l�wF�o�b'*~�Z?D
$@�!������pj'B��@�Pt�)Nta6�^�'fzЇ�Ե'�d�N{�hǲ���gv��GHeN����xI]΋���G�T�㫁ӣI3�l�³:'):�cK�`���^(��\��������ω����ir�<�fN$��ŭ
z�,$QKl3J��QwV(�
��`�d;d��7��%��)U������#�7�n�s��<J������4�nf3q�;\`���s�9��� �hRY<�����lR���0��w�x�Z/��8��Lb*�R5�P�U����W}6��Z��bE��K�X�s��r7�M`���.��ܐ�,�7�m�~���DKn��Cf��u�F+�v�\�����2�!��o�o��Ъ��K�b�Kh�C�����N�kUE�	ļ�m��;��gW��
=8�!� i����Y��!�*I_?�U[�\p�S��	�ހB�n��^�5u=R[�M:�C�y�[E#D����N�Q �v&-�
X뒷��Q�F�l��@�v~�a)�/F�1���0�Kڋ'�M�@�	����!��rn�8$dTD�ה���<��]��K:8�RZ�/�͘��m5w�8��{K 0����3�p6�	��;< ۠�V�	M��Q8�%�-�+�0�����UжgfE?H����(����`��H��
w'}�]|��7���$<���#�BGy�����]��G���:�M�Ӟ�/e@��E?I7J	��4��.��0�mB�8X����cب�����_�s�A�?$���7`f�(*���}���^V�DcD�G�1h1�M2�p�]��
m������XL�*:�D�������Y��|?q�ldKQ�a90��Dȷ��k���'�3��*��p���6�å��O��(������m�06G���4�fn�7@�}�rA���(�\���_a��l�eF3_AY�4}AC�/�8�)���9���6�x��6��єa���Bѫl��d�f�A*�F��>���R=
/f�zkg͢��޼{�[��zNx! G��:OX�h&��#:�^�R+@�o~	�?}{@�E���j���K�����#J�ӱ}	�^�^fB�+G%�0��k얗e��3��R�=�� g�0�~����	�=���j*m&���n����ƪ�P!Cq��L��*�!����p6�@S��&���q�3^"�XB�¤�J�|��Ҵ�)ΚۂXm�$v*���-�}�d�w� uް�
*S@��!-!irH]�iA�o��C;J2���%a��v
��(iC�
�7����F���i��2�Gl۬��Zx�U5�'�	��>�np*O.nj&�z�,�o���C ��=M�؏%xY��ׇܛ�v2g�wT��}�����ާQ�8[<W3mgQ�P~�s�l����u��N���|�L��#��IF�T��r6��W��Z٧/�k�����D�5'�ۆ��R�c`ҸY�Ffh!=΃�*��z�;8��QL�d���k_F)`���a/�P:�X�XΓ�m\$�J���mB`��iő�;D,}%>�>�0F��H��|r�'�2��$8:y`�6��L>��g6<��7�ܹ�E���w��Jx6�I!��i�9N�e�Nq1��מ&?��C2C1�D �������3�h��/WN��S��Ge�������
eǟK!zkş�o�-�=a���ZnK!�
%�O&BV3p��ˮ)t:o���chBց�;�z]�~�	�i��� �<�{���"���(I��ѓ���f۫�[ųَ��.C�iݏϲ�oT���6�#L�q�?f��pd���F�It����b��H�[_[\]-�'��4��zUO�Z��v�A��o\O{���y����)G���{��@U�#��H��Q~��Q;[6����h���Tj.�[te�&2&��&��..�7�~���S����0<�؈-��YR̈́�>.�2��3hcW�~�^}y����&��J®�?\��0��㷱�ԡ �%]�K�[�����ܹ���G�~�f��b����D؆��^X�PR��K��.D�.娖C٣�1����J�}o�By��Z����Y��R��������H�5��#�%�yZu�8C3���*Jk���*�i�f8G$�{z4!�7�_���g�th�6s0= 2��-���dEY� ���gpZ�(��ec�1�y���:��z�֐�x�gp�ms�X6�L�2e���%p��5C{Z㜯����ҫ���W��v������ڑ�x����K�d�{�.�H�cnC.Q���A2�))�e��hkg����:;Rdv�T@PB�B�G��'�&���cxف��,2���0X�qШ9t��+G��\�~e�\�Y0ZP&VZkܑ�C;�*.O��V�g:!����d�Lx1�q��@�*6��)>X�A��)Þ5�� 5�J� �SH⭧9����MB��,�yxz�_AJ�Q�ea�.��u���|�欍��t�2���}�۶v�<A J߰$Lo�R�P��"UA���ÜK�����@��lx�����v�<>
��7)��2�$�VP�2Z/'�5���e�֛�Aa�Q�h�h�5F������M�Ͳ�9	�A�N�/B���HV�����._f��?��I`���0Ap�+؆�e�A�Y��r�Ow"�&�SY��까t�v7Q�Cv�n��>k1��9�S��
/kw��#����\3���(��-Ê��a�&��!���u�����͟�Z��˓�h��:dÖ��RY��2�e�zr�}HqC�k��[��9�d�8�A�b�m��5�SnU�Y��HlY��O��T���J�&|R��ݎ�����f~bh�]������fRJ�^xQ�ȧ�$�-
���:6r��EfEɔ�E����P��F��p)�(.�l������N�@rG\%�hYƐ�dT��OV���hX�՟?67�\ B��^��~j����Y�	��qS�8И�?��E� ��b
*�dx�Z����J���t��U��?�N���ƥ] ~R����1e c}�%T��_2��9w�ˎ2�x�
7��@��r�9�(���X�46��C��R���.ax�b���k���#y�=p*�穳���ؙ6�N��`\��,;SFP��S45��6�2�� �OO��3��Qe���ZŤIyڲ&<��ׄw�v���[�}'n���掁�p[�\(ƌ���	�L�,�&q�j:L���Q��p�G��p��K��/��m�ZY��������, �6W�&��5<��ģ=F���t���!]}����Ѻ®�k�p	�l�#]�M�߃y���zXɭ�U ����tOE	&�}M�nK?%�}h+�UОJ	�8��
��Y�,�:{�r�E$x�f�m,�1�i
a�W��(�o�s�V�ؗ���6Enb��Y�'����ۻ��H!e{��c]l��d.���l��.�٪��&��+����|�w�
`�c=h�|���5	�9?�^��B]����:��:]6h����D��l�����_='���Ljʘ�.��|U��pp�%����Өg����T<i�J�V���;�s=mZ|)��찻�؇�>A�`�O7�g��7BŤ1�,�Ɓ�|�Fd �� ���۲a	y��g5��ډhQ�̺d�� �f�F��_�5���X/�47��hQ�����4��-p�˱��6�kr��z�N�G��4!�ђv�mF36����8���z}��Q+�	�� ��R���b0�!�=��l��{b�ԩ���}bמ�N~�&'�6��?t�=l"ܞ�ձ0��2Jf�i�zt��n]�!�H"6����B�Q�pp0d8����w#|��$L
�����
�4�F�� V�r��Nm,�$յ_�bWb�X�FF{�A;��[��Ɍ�
�c���� ���k���O��]��-`����P�b�^;>�$�0I���ă�"���xl�D��.���x���3@���(���}�ɽݭ��N�Cͪ4J&h��&xi���m�\�̞"�^�M��[t�$�0�˿�7佩��[n��u��o��}�����%��P��J�mwȎ���K��]�T��p���K����<�<�11�!Ĵ��Y�	
F�eJ�@>F/B2��B)1��穸z�N�ywy��FHc�`�AնfQN�Y���+B�l<�3�&T@9��)�̂�VS'+R�����Q��=�BQI��2c��D���+���܈� ����v3�e�|"��;N'����?���v�W��r�+�ǟ��M�y�9{ίzfw/X>IV�]�3��+%�@�����.0��W����vA���u}J/�X��B�n{�yK����*��p�U�d��§H����u�TF����ߔ�N���1oN�5�CǨK���6`\�����B��,�|���<��v2,�F!Op�?���@��@�E<'9b+���
�h������N�~�
敿����!���*9�� $�:=�N�b	�ș�ɘ�ɖ$
+��	F��pm�XG�� L�-W�"�g^P�ˬB�_Ǽ �����+���3�ǡg,�.��8m�ٴ�u��K�xlGp6�HEW����[�3�b�F���d��oUd��}j*�''��|��y�>�t��o���g���g�s5���Z�:�*k�i��i#��n��ke�e��'��_=C*
S���
Q�;���~I�\FM�7(*BHь���$Z�gXpQ?ؖgK T΅����%��'�7�~�Y��Õ��Q��{��������4�y��̻���h��7�L�)$�̷Μd�Z�>\ao���W�g:gww۰��qcr��F�H�J��<_��Z'^�׻:3��0C�6�c{�qooT1/]�ő��W݌�zP��j](tK
3q\��Upb*E�ֹ�7S���`��\�ѽ�<��ukDFR,53����ՙs�Ef4��m�dE�wG6��r�-M�9�s�)�G�e���29�=�*��UW�9���i�P&�?�X�z�s9�ӧ&��&�;��;m�����2 �Pۧ#�eFٚ�,xa���ٓ��-�Sh�aN>f-��&�m	cW�PxY)Xm_Jt͞9q]VӉD��h��GX��|%=��Zfj��\�H�Q��hT�˨#ˈ,�L��U�L�&��z�E��R>{�O1fN�� g|�`�q�wx�'q~Fݘ�e ��{ne��ֵafDdo,�<����/\a����KS�����0��x�}nR��i��J��3��?|�N�Y �PV��H��e�AGu2�� ������P�ԏo� �������qұ�5o!�\���fD��#�:���}a�is|
+��5���;�}atGN��:�x�T��WS�4@��1���Np���uYё�xK5��\����p�R�"���Չa/g��̂\�@ͱ�N#�?�)�(��u,'����I�F�%�4袑Y����T��LOQ���r(����\��i�Α��/�?V�)�Vu��E']�J��QVU{x��GD��x%�?\-���ֲ.�_�<��ˊKC#���K�Lw�������tSJ�.��㍾M��O�Y$8���B��?;Vv㔻�Lt���i��b~ݳ�f�ɷ�e�߂n$p��ش^*�����cU����N���� XP����Ԇ��:E8�ưe��M/^ ����������_A�g/��S����fYR	�2S8wƇ�l�����"sh3�WD�[�o�Ew���Y�g�V��M�_ǽ��$$\��Z��8�[�@�{	u���J�=���3E�B�+���Xru�X
����$McR��#�ɳ�ަ3��k�|\n��1�^P�$#��>���|Ԋ�$Fo{r..4Y�G��2��2�;�;���	����i�!|�z��gs�E3��]�oKV�����y�8R2q��x �â{�W��E����l���ө��;��h)Dt� 6�<����ʚ������Fϐ����1bH��T mB }�1��;ځ�qQ�	IQ�~�M���l��ɑN�8Z��9�#A�~��s�L��oN�t�E{��!�|�`\0;����MO�M2��K�yP*>Q������= �
�RwEF�೭ͬ�A�ᢅ�S������z�F�Il$�>a�Ȳ�7�0~̦�C!���K���q`@�Q5����2���Csf�1\�0ɚ��,��r���۷yk̋:V��-*V�H)2M�O�^V��h+`���K��3�Yu�T>r���\��W1��X��/���Ta*�c�0��d�A�������w�>uk�&�]e+S�f^ ��^�6g���t۹�B^��A��[��ӓ�8�2d���2�$�����L�O�c��i��t��K:]���l�Ң�FڳIS�x��B7��T��z�b�q��>"q���׵�9�����j�Tcqwp�hRbǾg��o�!)dt�̍7��]1��`��ޯ��� Z�o|��0;π>�d]%i�ɚ����Mj05Z�\�:�	4C$v��5��Y>Q�~�1`�K�m�-�a��Z��NR�	v&/&O��HG���^#\�W��R��QyQ-�m%�{nv^�ӌ!�@�@��IW]����}��f����=��ĥRx�t��;�@�]yĀ�r�fP���8w�=k<��#�U�G����Z�-	�d1�3��s�E|�����5�/ݦ���9{! r-�5�T���΋���K}�����'M��5��'��`�z�jP�eщ;��ӁC�	��,2����eϙK:�ة�������g���>�W��nX��dKg��B�f�z}ר����15
t��7Sr�g����)���Ӳ��ʂ!�(����4�k?���ߣ���n�Ѫ7[��aw������Xzj9�����Äoq�-H��es>�\����Q�k{s+C-yJb󣂅!c�8�AȮ��&P��%�:?`><�ù�qz��gȩ��e̊��v��oT��ƍ�=�"x��@d�k��Η�-���TX���Y�Yr�
���]�3
}�K��;7����[45���;�)��܌1f?��4t�,����d�I/��l��@�b�D�r�� [����a�&�p���K��ղ�o��K���Ù��Ȅ1���L��������I����m�kp���C�h���Vq2���?r���j�:�O�q�����uB$\>���d'�.��TZ�Zk�Ҕ��q���|���&V^���skY�/��uʙs$�az��{�_���0���fʴi��14 �&�]>�apCCwt�z�'�֒'P>6�����&��F���Dp�s��,E^�X_ r2i)�2�ltGF���u����˧6s%�)0[��Mq�?@ysr�Q��=}P�9�t�e0�/�e�ho��K