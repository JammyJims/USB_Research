XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#==��2����f�r���"��>�o�����1�Q��A��"���e0��#�5a�3��RD�S�
�7��X�ګr:�,s/�Ç�m��yw�»��g�j>��7��M��/�恴2�c�%W�G���+�%`,	���եī��u�!X������h�#����\#T?o��ظ�k���b�����.�#Y�]�����	�G�G����H���J"Ժ�n\��B�W ���ո|��͂��-�#'�z�pj�gw�F����-P%=��b��3�g�T�,R�b]=k:�aƏ3~0�@p���� $��^���$�U������� S�w�L����� (�N���4��!���0l�f���zJʒo�Ř�+.�q�u�����ea��\�u"��Bʬ���=H���5b�����IvK�Q���P��\16�m-�>D�,��+\����żu�F���I�LT�L+pjw�5��w[g {ٍVR
�Ϙ_z�
14��=�Um��MvE�/��j�X(N�`3,3F�����'����BI9\	�}� Y�&�(��G(<|rW&Y�S�{�1[�~��:2�&9O�鉼�+` jkI�G͛�S��C�x����:����ֆ
^Һ�Vh�Yǀ8�;�F�3��
8���^�=�Kt[�uD�z%E��=�� %��cbAh�	� �G�VѤ�#B��N�eZHY7�
���7@0h�V�)GF�!�b�I�l����Lh�Ϻ$���xXlxVHYEB    49af     c70�W)��� 6
�:���^qco�]��'����T�Fz;�p*Co���ZA�.́BWM�+y�C�q�ղ��:�D	5��Kj:�!�IU.ۨ�b7�F�g[-]?)B1��6c�*��o(
&���gD��<�31D-i��{(���@�A�Y��27�ʷ�R�͘��i��:�7-�T�e�HW�w��C)X�h�GG��|.)����f=	z��#6\ټFص'��:*Bw��p���v��A#�A���_�C^�x��Gq��Ͻ4WX���0�
'�'n��~���A0�XY8���EK&�@=�!�_��9!��N�Χ?��[߭�"sھb0�/ ����G_pI���e��Mʘ�bv�5o��l2����FҠ���\އHp�p/����k�"�۲��'��@���@��UP .Q8�G .�:�41��R��wy"�Ip���K{
G�ߙ��2m�BǺLx}�-�$�A�o�r�\�Ȣ�b�4p0�����o��W�|�5�3 M����=`!�9��-i�R�� ���|��|e����c�Jj���n�S���OU��ʞ�����S���`�a�
�G��A߫�Ѿ�ubT�m���Z����Bo��x�
CT��؃ϬEpg���gb����o�5�͒(���q:Lѧr��K"�ߤz�խO��Z��ƦO�l�+.`��؋X�oEx+�Q�:࡬`��� Dx\�i�a����G�cɽ8����wSC)�.Y�Jk}�_
�M��|��$?�+��=>Y�C��Z���x�9痆�")����y�XE#��}RȨ4a핲�sX�?��8���ïD�HЮ�@�n�k�#�1�9Ϻy�Pc ��>=8�D?a��I�7�����6��E;�GF�[���lS��	Q�>)������w�6��.����}��cˁ��-b*���R�:��e�*!כ�M 9�x�\쵡b �-�NTȐbv�ǑT�o�]Y��X<��o.$���7�m7�ޗ�;��1㭲`���p�`�	
6z�X�A%r��.>�)�ж�Z��88����Vv�Wm�*��O[A5BG9˥DNf+��S�
~.W�M&��r7��y��M��R������5�1TK�5 ��9�3ߩ|�,�U�98f�� ��2�n6�e��sv��|������]�o~;I��[W��V�2��,�ԨJT�g�b�눈i`���"�]w8�/���N��Le��	7V�����/%�
���p�<Kό��E�Z_�����)+���}'�A����*��U�N��A��AA��W����vW�o��U��ʪ��@�ÆA3`�ſ��V���4"��1	q�u#4���A|;g�w��rlO&�U ��G��nLIZ��/�/L�x��G�xN��m�'�:id�Iܿbqߞ��CqsP�c���T����'m��#
����_s@��z�Q�u����m���@�`����[�ݲ�����"��x��q\^evEB��7z@RB��k�s�_ՅG��H"i������}�~,^!�z]�?��8�)B��I&�<���8�A���P��l�KF���O�����N�����-!�;�3c��{Q��`{�'��[�d�a9�$�G�H`,O.�%Q�
�������v���@'�K����:x���y�p��Z� a��[�ﾈ����e�D��s@2f����qB;�G��Υ��D��L�&��l�^�#�0{�1����6s9k�~S_�Q_�T��e!c:
��(����3(���3�[�]�ڧ�ʮ��<��۷���n	��/��dFp�����u�n��K-��h�;�wg>֧�����cfCy�Z-��#�-V��:S\T/����'�$���KNH<y�%-��O3��C��ln�-����`��gl1��Ռ����58��*���U�G
ј��?qY�m�L�,��2M�
k��1����)"T���Yz��,ya���Jn�#�k����^�����C�:�mO�c|���>6��(��EI���oG�U���˱�/a�vI&�ʥ5#R�ח!|���-�7��-۩�)�����c�N�Z��(���Y.�a�}<�\<C�ܬ���47��i��E��E���1	�h���&|]�(
�#S�
"�}��_IT�1(?=r�<���}��":���OYZ�[di)u♩�ʊ�;`����2��*�(�vl��5/�T�D�H�������h��(�6��
Jrl�@7g��_�!�b��n_Q�X��6@d�7q�é�&b�v!��!�D���V�ݕ��}~�fV������nϚ���
��t[G�����P![�����i_�;��+�S�M��d�%҆ƌ�$l}ē�� %8V+F�5"�"�[f<����7��VϲG^h�P�s�Yl����V����|z�wb�;���L� z�Q� ����=s����:{�R���~���f��w��4�Ov~�̜7�ض��YB�+($~�S1�ymOT]?�R� �����bc�`»�I�r����r���M'��E�5`���6,��2��.E\U�C%��c_�j����t�"`��`�`���id��m��F4�;���	�I@|$�0���Læ���w��B�l��{t-J�u�O�߅��ݹ�N���f}�>rc��+���^�St��	��u�^�J�qD�-��te�Ǽ��@9 ����G���qP��C�F����Y!#� ��0�/t�{�
5k�s�\�'���������]�Q�H�[����n|��`ð�8{���~Ł̡�tw���."���q���ȝ����si��Ĵ"�:������~ᓹ=ބ3��Y"��I0�����1v�`��R��EiS������.��2�:l�f;�9O�M�6��*�hi.��2�R�(������q��<�fꨪ��a虧kX�F��2`^ц��V��A�ŀhKe�+�+��k �Q�Pt��l��*j��=����|�ѧ:�ļܝ���Ե�ĳ����$�]K�L��u��xcO��s�a�+�Q�?�������l����o֟��ڲNc�d�TNB��C#_Nu���?"��#�.��DW.ټ�?y���Bxk���*~�j:�