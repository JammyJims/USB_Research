XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G�Qu�
�ػݙ��2�r�t���,z;���Gr��_3�9�z<���:aE���Z�ט���OE��ܞx�(I�!_8�,�󃆼�"��UA.n��m�&�7����n�h���>���B�L�%dfέ[��R�z�-A���*���$9j�_���} }�EW�&���J���᪉���#!z��2Xț�\'qȖ*��7�N-i"c8��%W� w�%%�Z+ge%A@�O٤E֝a+X��y#B���كO�9��lX���\rr�1�v�� ݼ^�ԏk�)�	�B&���7y3��j{��fMHE<�y3�Ed_?C�Q�BZ����t����9�6ro�pmB%����_�N���F2�8-�xC�r�y�G6��?6���j8��Xv���H���up��_}�;@(��z\�H�2����R�g����:���c��h".C��wD�P��������T���� S.W���nx�}[3cd���v�Ɓ� ���ɵAi4�$��bq�C�UB?I_@ꡧ+�D/?�73-�&��RWoH���lkr&n��'�x���
r �%"�ޫq\�jV�;q8M�+�#��ܺ�����gݓ�"*X~�IC��J~v/3o =�曙�}e��2k�=��Q:Tl~��x��d��>�&s2ͬ�0�è�!v�Fg�2��ȵ5�iy��t���p�vpg46���郵���΂lU� ��߀Apw��X��u�XCh�&�0TLd���Q�,փ�/�U3XlxVHYEB    10e1     740�*��P�6������Ay�|S�Mv���$�z�m�f���x����W�����A��s,�m�A�p������A����$v�|A_;\�AY���^D��V�hr��JA�Y�ő9����?��d_q�w`��pYĸ���s�n4����*����Қ&j�ݵ�M�@e1���Α/��iŭB���ki�����#Q	`(��u�s +b���ҫl��n:m̶���j^=���C%��A��3������k�����	9�j}큅����[�ܜhIɚ�)f���-��R���PF��魶�/�Qu"�Ahyw#=���P-�3{���>>�y���x����4LWbL�k�F�� 
G�������p˜&)�k��lJT�]��ېW-��
an�8i��ù��͊�"���I
Z�>�liYSX�r1�O�yD��>H��moi��+6[	d%�ot�kl"����]�!6�k�M�ݙ�S��������8xN��]E��Z�c�Il��3�h��L����0�Q㨬Fq��I��[�G<.H��;EF�Re֌��c5qI��|4X��\y����UZc�\�N�;�g=
�clV�����B�:1M��/�am��Z�n�T(J܅V�,�ӏrA�y�hm���|6�{�TJ���Tq����?��긓���Q=@#`�3�/s��[����H��&2�༟��	�_ �*�0���HE��+ǬE�>�/�B�w�W�6�f�>�վ$�h O�t�z�-�]����u'����@ �� �?��'��x�q{�/�b?)�рXɐ�T�k&��ک���-�c7F�a�4)�h��~��v�3p��!򓽜��J_^ xC��ڮ�g�3��,-V����^!:�L��%�R����ks�H����|�.y"v%
�Ac"�q���G!�����xa��<�j"rʋ3�C�#���2�#�.��i/c܊}jn4��׹7�RL��4쩢lݠ����9��S���>��;�uP�%������
�
$;��ՌyE�j��@"�]�a��������g�˯��wZ:m� T��T��>�C�Vb�Ҡ����f�q�r5-�Y��������������!�c!�v4�,��cQ&FF�Vy��6�0��E=�J��h�]�Vx"6u\Ԭ	�.�8�]�����F��G�k�͝���Y�0
�%z��4rg@*i����w�Ё���Z#�6Bǆ��K����P���	s�DL����t"�a����.�$x�sL !���g�Y?m�bN�9�3ؐI�RH�?�G/w�CH}0XnA[I"v��X\n}sI"?�%x̻�-`�' f7�x���\�L��v1x^k��"I���O�&����B������)�62}I�+�4<(I�_�Դd�q��^�Hn"��2!(�mm��8]���f�!���',��oL��\'E?�f�h�(�_:�Ӗ�ڣ�2�G�F�Y���9�06C�għ`��s�0��3���]���
�g�^OVt�]�׃�S�#j�Y6�y��ɭs"6"cn�:d���Q�ZZ����{�mBe�:��D#��|jU��J�m7��c��Ş�U��69�s�ܦR ��i��9��r'~���V`w���m-��������C0�iQ��lG8k&I>z|��,N�Avsv|�I���6��xՊ�,��o�.���3]z5	��O]	�N�ߙ��g�)$��vז$du���Mpڂ�A�/v�0X֌"��&��N���Ày*����;�0���W������ )$w�
[�Ay�� 5�i����lGƥ��=�����4`lF�Q�4{�=LN|��O�����ɬ�U���/^G_,o