XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l7�CI���F�
G6���s{��ˏ{�S�I�h K�*xބ*�)܊8��O���?.�>C�Hx��j�a��j��\Q�W��t�iߖ} �C����V�C�9^�4L6�/LuiH$Y�P]���z�q��"A�<��]-&�f����T�RV9�5���ly3t���!ʗ,��ld��PO��Rw$���5g��b�5+�i�X*�<�2��c�v"�	��z�.�k -� �l%�aɍ�j8#�9�'�i0�3��5Aɀ�#`�?<�A[ׄ���=@���-�6�.�?��1���0c��9�x����PGSh�A��9�X��
�q 9�^w�D�8x	��1�-���VV�����O�A~K���3�
�g7��O6�Zk�y	 ��]Q���'����K��p�f <�J�q�n�ȨA1J�T
�/q��%�	R<4F�Z��|�ܶ��꟪��쉭z�'U�n8ƿ�eg`�n4T�t��̊���b�LA�������8W��'��O<f�6��&�\RR"�o�g�$�$��fK��#���/��h_�`�Er��&��Mh�91]��6Aࡁ5Q�_��qg{"�^e����ǥ���	1˓?B¤����w�#>��v��}7�H�ϝB��Am�I����j/D�3���!Ǆ`��x�M�sX�H��:u��>��E�J݂L6����N�v
� �2V?V�__(j���H7���"Z!�B5�%���4��J�Y��U���7�"N0�'��XlxVHYEB    49e9    12f0;T\��3�E?$d��Q�L1�{,�_EE�]Z��C��ad�`���ZG�͐��H*�NGl�ґ'��<�#��sJ�؃J�%�n�/)RS�.ݻ����MU�9����n
unE�P�d2[� ʒ9���X�i��T0x7?O,��H6b�]9���=����&�|L�BsKъz��H� eS|Ӝ��JAl7�����x�)A�*��h� ���3Ci3n��Lev��͗Q�(�R����e$B)���
��b�����T���`8h���w��	 ����Ww�Eit��s+]��dÃhiܾ��IK���'��ӓo��=I��k9�����tq��K�.�n@ϩ�W�%f�������P"�� �5ٵ�.�L�<�2.�U��M���@_��1%rs�[F��	�"K�ҮIYC��Ӗ<T��`�Xod��g_E�T�F��ƤPYA�i�M~0���+n\&/s��rr�¶�*a� y�Ky���ac�!�u�����U�kyQ�T����+c�ЭRe�i蜕�&��98�=��k�e[ar�ĭm� �]
��	��s:��ʽ��#9M�^!��\=v�#>W
�;�V�Ln��TS2���r�
����*<��G��ˍ7ߌ�eNFl$4F T��lU���$�y�TV5�O"������'.��t�z�[�޵Isl�D��/¾6	����|#��-;F��7<�τ,?��_�����{���g@a�zTL��R���u�m���,Ē� 8��pP͓Tq�fB{�Tx������_ܟ�cF޸��[K�S�p��e�|^E	�$�]���^b��9]g�PV�`_`��1��*���o��B��} �1_c�FY�����t}q�2�����_>�2X��_��51��"�t�9��m��r��1H2gMGz���u�ۓ�Ч�M�3����E*}x����T���ʯ˖�O%���ӹ��H%^�pt���ޣ���
2�P6�)` �z�C�ޟ��!��!��"߹	T�G !�^7<8�I�ӊK� ٪Ƙ��2y&�gE?4�����Y��)k9�L�G�/T¦�}H;d��I�`���{��uCe�4��x3�a|��i��r�Ս~"�h�X�i(m�Mo�Ji/д��KK��\f6�s�5�R����%��[��7�?�E�X����,�!*!�E�1i���s�(Uڲ������Mp�
11�����Nk��h&���(y���S���/OK�����_���BE��cl�f�2�q6�g�yVvs�$��1�\`����~�ݠ��`���j�;Á7ߋ�
4�p4�'0e�g! �@��s/dWO�b�6�����U#{H`n�\w(�Į��.JX}�����:��N���]�,*���;�9��-WU���?�vw�٢�(���}��$2�:�����}���^3^)p�5����q��>�-�Q�rP5 )�T� s^�[ld$V�#&-BA��`6�8�A};T�a������xG�s��?�wcH���  ����9f�_���T􈚀YC2�"�4<��mb3�_���[W�c}9���r7)~�$o=9̺%��@�}W��d�M�S㢄x����jI��-�\���;�����f�ϱ�^�.Ƭ���|Z��>u���~�j24s�3��-�'��f���ɪ���$����8�.�_��G���m@WF�c paL���nD�K��ڪ�V(W����uc�i����8�1��(��E�&�����U�n�@�/�@.��n5-ߎ�4���׍��yA�x�sT��rJ���+EqT}[�I�tGE�m]�m�劀��̣Yi��=�ǻ`:~��z��9�
>�������ʾE ��e�c�яp�|eO��9�k+J�A&%�g3�M��&Nu�QH�l�Xԅ��  Ra��P]'򈤸����m����r����O��4�<X���"����y���S��㘭��t�3'�HP~|�tJ�ŵ�5$�T��A K8r�6zme'�C���s1&R�	�rϧx��v��4��fz�^#SJѭ.h�y=��ҧ�(���͖z�g������Y���<Ч�ّ]��p�	><ӎ�:<k(r��ˡ#�����좡�;��,Cʚm�ǭ��#v=�^Y
�6/�w�A2���b��\Z!tU�K����#n��f����tQD^�c��Ǆ��>�hM��|��F+J��nB��dz����+���X����,*�����@�|��2��_�� �&��-X�'aY��/P�_�`�5�WY�lTo ���v����&�5C���d�Nq4��p[����bL�O��l�Zvul5�u7�\��^���0)_����d(����q+4��D8�߂�@k�;k~��D�d���+�M��� !����r���2ڝ�5�T�
U��9'6�A�0�Nً���]O��L�j[�$DL�3���_��$9`��fˮ�&����%��!��U�s�O�=E�i4(���c�Ap�MC�1
�ڴ�_�&sLh�%���D�!��I=Q�;	p��x��w�?P@1�Q�^l
��̤s ��o���w��sUԘT����|[�b�A9x�ԠH���s��Z�U{	�n;�{�>4��xSA�&w)�i ��@{+(�ۂ*P�X�߼�i�U��RX���$D ����*7����>��Hf��R�3�=�[�oZ�taЬ ��TSj�Ҟ�Э� p���-�)^;��8a�fT�3#�W�u���;�h�n�xQ�0ySy��=9jX�Hdw���{��* P���X��95�ֶ��ʰ*�:�?�2`U���av��I�ݓ>����e���GGS�N;�h%�-�����������S:���OLƵ-��9�*�%��{��@�7�uc�ש���/�
:*�0�rPm�e'Zf��|^�<1�����S_�L�hBPVR�M .��"X�Ս�ޡ7jr�r��@B�����f�����!!	�#��L����>7����ԯ4�`�p0�~"�\s��a%��z?o[�A�e�áL���0A�W|1YR��AO�!Ue���(�!/O�n��V���ؕ���l^������������o���V��Ƀ�'�ԫC�:B�n�3�I�(܃�E]�G'���.��a�R= $�SW���:�9��˃i/�Ό���T�.�dd���������CF�(�~b�-���a-t��7�G�������X3���ߗ�z'E0?H/�FW߄�t�8r���o���d,I0��@W�8�V���	��������dq/��a��~J���,g�o���4�֌<j��6Q�I=+��}�B<�B�r$[�Z`�<`��l�vh��p�}��<�'Us��\�y߰�x!J&�\��7��Ĝ��b�O�?��@�5�K:�p}x�t��4~��0>�7ޝ6���et�!�;�cŜz�B�C�F%�fS���5���5���[�Z���t6��]hQGd4�0^��jWQ��9�Tz�U�d\W*X�8@X��|w�%���܊�C��t5�9����o���ի��G����.��i�Pz]�kC�d8�������Bɐ9A9�W#3x��}59��$���c1!��-���`6^f����QD�A蜯g�*�r��쑘ls�����0�`N���O�ѧy�|P|���`�e���$�)�ra�D��W�E���rgKu�ߦ��.�q��z���Oĩ᫮�i-zMv}*�_7m���,�5���2SsE�n�JO9V�U�����Xm��0n �.��G:p�aꉇ�9�rل�HArL���~�|H���G�u8�7�0W��[������ٕ��^pf��	�E�F���R$��˟Bsn�����X�3��������S��e"#(�\�F4=�'�Z�Ӡ*u7��3;ȧ�K]�_�)V��h��z�3X�F,5�?��^���T<�*³��(��&Qĭ>v�f�npUB���T���<8+?����S�#�5FcЎ6�CaįX)e!Y��sm�I�]��/�f��̥^��N�{�9���yL]8�5�5��ya�L2��ҼF�:p�z7g�2Y;��W��描]7�4n�z^�U6JV�(%�y�eu��e��R/����V冀�#ӯ����<H�T�Fhn�����*�ʥ=�(�5YX?F(�ۇ�^h��ɶX��ceo���f��^:�+��̜c��-��[�D|�=���ہᶤ6�dZ�wު��Q�;gwF��T��L�T&�̪� b�S]��u�)	a���`�f�`#))E�R��H�/ we(nO%[��J��� ���&!��*y��\��&L��2Rd�15��.,�5�=�/�������Ѧ�??
Z+�團���w{�ǵ�|J��ޠ�(ɛ�t9eg�+�!��!h\*���7��l��7F��Qc�#p�b��&|`Ekl#w`��`�9X�m`�c������Xb�j�>��xYmQ ǀ� 5�6�`Ѯ���\E^bgu�J�ػ2�Q�����K�22��'�*.�np�<���brU�VZ=����lkD��<hI٘d���@��K��(Ww����"�0���J�Bn[{���([�s*�|�Hy��=�����������[+Yj��>���0=W`�p
���8��]K�e�aó��(�s�y�M�%A�꭯���g��x�5=�ؚ�6�l��@}Y����	�g!��1����Xm��K�%;�d�RW��qQ�k:�I-