XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#�Ku��m[��)�Ff���!�M�����;��eҔ�`�:�[3Q�c���&����X���I5��^T�E��f�YM����6�!Mw�V�����f�q��
��-Ps�e�ō�J[w'\.��4��A��Ƴ�(I�i�mCѦ���FȻ������2��;`g0��hU�j���\��F�S�T���,Uʓ$."7���I��� H��*�t�h��$L6#'���Z��mɈ6�)��W�`31<�V?��I�?�It���)��ֹ�	���Q�G?�Ğ��]���ˌ�*���0:��U��tJ	Ix�h�b%�r����N1���j�T]�p��]k5�V7�Aĩ����7o�	��,Y1�� �Us��H=�%� ;�7O��-0�k9��U�5��m��v��P�����m�w�ĺeoLi0�.�M�!FF%����(L�i����&<g��H$����:@O��7�R�-<��|��]>��s�RhA�-��ǫ�T6�5#��LL�H���Ԓv���c�r<���.��>�"⇪��_Ӽؙ�ěrF����%@���5����و���Թ�����0nZ��;�;�꺊���[�� �dA�482�<�
�t�G�[��as�y�o�z�"B�&�ϩ��^�B.��W�Ps=������f���՛ǆ�hB2�v�,��A��{�
|��I�O/ˢ~�E��p4d;�{fQv�ub,C���ΞJ`����~�m������*u�<�fXlxVHYEB    91d6    1c20ƺhW�]�h�$�e1H&���[�R.H������bx;6��/�%�ŲگI�r�*apk��g˝�.����1��,^#m�����o+����l^�팩�tʳ48o�lci����������5'%5���N�	D��Y��$�yO_�nT�d7G��P�RBf%%�{p����A
����س'��K;3BQA#����q���9]�[�./�9r��A��[C���[�yϝ�v�r����D �����/#�:��r�*�#T�0����[��[�d(|�����dWI�\�M��S<� �t7	e0���v���&�MZz7h	>�b2�^2����3���	ԅ�2P�#_l�]�
{�B���$<�Y��]T�h!S_���?/��._�t�m�ck޲@����=(a!z���o��fsaL�g��0�2Q>�X� ��3L؉_�Ž�8:H�X��l�C�~�I�1_�2��
�A9���e�)�f2���_�z��W�d�<�0`Wy�D�U�O����ۀ ol������׸��i#�tQ��/'��7��Y���m�R�ja�Q`A��+mnL�}M�0���(��U����O"�s?�Ea��*��:�1�2��Wd�8(3m6����^�)�گ��KK+�@2��	��1yfG���x�6N��%ݥ�;��iԼ�� V׽�A��Y�|���Sz����c!߬*��e�9� �bi"U����U,S�G=@\j` ��ݫgވ�A�6�; 5�jڇ��G�BV|�/�K�E:S�umD��1N`r�/���	J�#�r���a����]Ÿ�)�R�Z���$������$�@��P9��G4��Xlb �*Z�Y��-^��I���0����)}d����鿅��X.��K������c���XHհ�4Զ<=9'��5?K/j�I.0;�A��8��vN�ՂI�Pq76BiQ}�����>�YD}@z/��:�����`��i�+qP�B�G�O.۵� ��7��sI^Q���>E��k�s��݇�_�tM�Q�_u�C�S��(�;Y�]���9�spp�=n�*�?.j�B7�;��	,�q�[�>����N�l$7k��P��A;S�m�����(r�>ޡu�1߈���A�Ȍ�Nl?��3r钬��'�N^d��V#a0�,��:D��i<�q��td���8��ު���v�U"���	n��w�p�GRy����
���e���U�/��$������\�Ts?�����8�݀"�_G.���T�:'�s��4�E�`���-z;�~��w� UHj�攆����O�R�uv��}��`�eFE�Ɲ�I3P� b�JΓl�n"�U�^�
���h���1e)H��׼�##����36RBv�sٱ�o�lm�S�΂�S��f�)��2\e��m	�횒�����.V�����}4=��4�p��6~�N��
�h��W��J�;75��y}ueXIe��p��a�M���6�bߐzi�v�H�G�O��j�SuXO�Or0��_��;j���&������;ܶl�yS�j���Lǝ�j��� W�im=�x�WPc	u���F�8�u�Ph~S��Xn�K"ׅ�='I�p�@��(�ч`S#=��M�ӦiG#�7�O��i0m �!���Z����j��]5�A�V��R Sm�}��<�����:۾����%��� C��6\�i����X��m�f�Ш�O�Ek)�r�[G��ȧ�mbx�ntGM���x��������z� P
��R�ژXwI�� ݥ߹�Zp7e-[�J	��4)Nnc����)��Jk���"u�u-=� ��7�RD֟䀇�	h�e�2fV�f�^p�)�P��v�2C���-B�2��q_h�/���
����,�ظ�n~G��nu=t������F��&e����^l�Z�?P
���2��4r ?<���=�]��88�:��S+}4�.�2J�o���x��\Vu�Z(�4���8 �e��E�%� p�U�v�P\s��)�`�g���%iP'M/�/�>���	Vf��u3^�����v T��D�Y����BA�B&و*�s�U�]���r���o�yW�A�ˎ`����46�MMO���u���=�.fH�P��@�jt4�4m��Q��/GfG�SP���t��0G.'&�I�a��:����%p�BX���6��m��!��'<+	��n�Ëw�B��`hz�:4@��rb!�u-&��e��[̔:�|W�M�ݍ`��?��i���l�M�	�I����	�S(��ū��֘mhLC(N��a�A��DPz#����8��u�0)��iU��ʂ�Y{Jߴ��r���8�W���5?����I�����b�TO�+���y�D���⇠�I�����у�/��X��7����]�'_��$˛�#p�
] m,���	�w��#t��\�&�+6�1L=��B������lk`���M[J�e�:-�(U�tS>���Ջ@������9P��S��3���z�������q���i��Ś��9Aa\	s�)��.;�r��^��m9��Pcs0.�$����^������S�gf�\.� S����@
6 �Z�h�&E��V�N}fLƳbWs�h%+��䯘��\HW�����(����8�������_�n�ô��4��i�9%��Ϫ^衧Iq�3;��!��3�W nW�*�i�����ѽ�?�l�aT�}e}� ��y���]5�i���n!^��K��s���3ƚOq�Qg��#�A�'aR'�w����M� ���A���%�)ƉV�N���T?��w�ǽ��n�T��ϔ������+��䍰�P�����܇rU���(̺�yF��b�u�ہ���RP�B�M;K�e\jJ��$�aeՀ[i=�f�ʱ�f�^��H�_r��7'�kEE=��z$� �{WR�R:>3TB�MT��o@��1QH�2��l_�X�}˶S��m�&0�qs$�%u�BGV�9����Ə����������ʮ����8!�U��̝��,�e�
4LJ��"Ć��$���#�t���b��]4�a?�����^��e�������2[����}?�$ш]�;GB�9i�qd�Ll�.�D]/�onK.���ڜ�Kb�{C�ƨI0�����ES�Dv�묒�ɢ���jZAU:�g̥?��i��d_��欥��]y�Z�J�:�.}������ �����t���æ�K����7��Nl�b)$r�t�7���G��ڲ����5}z<�B�$m�B�y"�v�����S�P*54�O�O�+�F�����Ex)_��F�kǎ�Qo�K����������Y���\�_��,l�0���3g9nG�LlI$�=m_9�FH�E�o�X$ȡ�`�6�#:M����`�r�����eh����Iq.4�Z�H=&scL���ccP�1�eJ�������_�V�21��ɚ��\�/)��q]6����0��fK�Yj��j��Z�A��e�iL9���d?�iЌQ|��o���W�����РڭE�J�o9z�폪���:0<7=��J�<��+vcS��?��B��z�1L<z}�)�]�'M���~�ǑS�bk�08/�%v#O7�Ϥd��)��΃����<r����y�O�F'Y	C�ʶK��f)lw!�t�Fw�<��Y5Ů�5i���y
�չF�\�E���m�Fx�ڥ/�w�nr
TV �}��7>�H|�H8b-ɸ������i�4�2��h�$V�@��u_��\�#F��ŉB�[�S��6��ʗ��؊�n_�%G������<\��9+�!�<Y�;XU8�2����L9�"%��s�Y��.�<����4�sJ�SHh��/&�cc�qmso��i�i��:}�(�>qG�c�l^��Uչ��UB����*܈�	�96)��J�Z�.����"�G�UB^�C�e�S�y�.�]�+�3Q�O���jl$�����{4ĎӦ,���R?� $Oe�Y�@���Gz{�H� a�<͕
Q��o����kb�x��AIԨIk�S�՚U��
Ykl$�m5�Ջ��r5�	��h���|C<6I�j���C1?/�	�ͼI�IJ��`Y�����7�j���u�cA�5ȼN�����K�sn��
+(����{�'B��:Mi�h_m���A؀)��v+�D7zܼ"E�T	u28`���T"�*�Mf��Y4=#�R�4ѫ��J�HB��LNa+��GL����Դ�C��[�2�J
]MlI��F�#p�n��;��8/q����o�ᙓ��|.��C��B�%��9������&��XH��m�}�D����%2uH!�4��0	��h D��5��k�x�9T���k��>���C�f�Y�bT��QSig1��k�E�R �ɐ6w���ȩ�A�e(���[>����^L�0PT�F$�"�}�Ty��9+)���!����?+�%]�Pޱ��F�\B;K�a\9t'0�^�&�`K>�l��k�c/ٻ2+WbC�bq�)?�z���=�׹�h��)�ҡ�ԕ��u/�B-���Aq��o����N�Ǿ��=�?���L����'��ȷ~�S:�����	������9�3����Е��H�O���Y��~��2�� p��uD%A��5H�)&'EfZ�H��Y��Q��f���}u����CxTs�.��ɛ }�bDkh�#�S����=魹>Ԍ�%8<����*c�,n�E]�q�ʌ�����C��1K���N��a����:�{�
6�⊟������C�+DT]ۑ�Ȇ�3n�E��6[d��eN_�y'�wAA��W�=,(�\T�75h�Գ-h?�m���f��Z��xPU�zYU�1m��Ȍ��Q�v��A�R/t�ϒ�J��V[�Kr������Y&�|bO�D��'�����+�E�6	������+]A@P�e����$ńgl.wV�$��V
a���D����/���D����LGD���IW��������[���"����c�
�O�ǧ?�V��=��SC��P5X��9Uk�:4��u��W�_��ϢF��@�W��E ���9�}���*�]��֡�0�$?s�xs�.ȓ������Us��#z5Q�o� ��Ç�XW+}e:$
��Y' xj,ض���IbFQM�-q�ؤ��(흥�SJ��$0-��C�ۙ/5$k�+�Q_�*�m�3�'BT�כ�1��a�C��PV�;��A>��p����-� �]x��TY�zt��qa$
�|�]��.G�cԮ):𲛜��q�p�?�t�F,�w���5U�$�4�*9yP5S�nY!��$Y�"Q�Y��޽�?Sh�aN��-Z�o�R���c�hIZ�Wa�Q�x 4���>���F���f���..�񯳱m����YS��dWU�� ��U�UPA��B�D'�ϒ�һk}������?��e��\��F�����M�<[sޚ���v�/z�P�|E$	��=#~��c��xgxf��$��2(�n�[*���#{+A|��>��q�)ё�|4}��� ��Kd��RCM��3.��q���!�C���;�������'P��n��H�d�*��Ɠͥ¨�aY�ب�B��e+͢�Hx������+��4���n^,�q�����nz��e���`���%Am]�h�+ڏ��ͣe:I�uz�C���>	 �GB��U��#/U봽 mԯ�茧���ڤb��'$Y\��?RAd��Y4�*U�7w6�
�Y��1��}�10��4 �$�2�A��񌲻�]��h����=���p,���mPf⑌_:k^��c��ɪd���X��j�K���gw��q�I �9��Me��
#M�3��$_X"������Ŀ���,+��k[�+5��>w�#�ʧ�dU����1(1��O8�(d�9�!���+3�[~�e�v��"��_�r�Zg4�\�����=M��7�`	�n���+-(����-p�5�c��#w���R�u��.A�i�����
����8l����PϢ���-.����@,��*O�s�T�ԕT���]��n��oLh��7mjUs`dA��N�XŜ�ͼ�d�.����=,�0�+3z��xn	Ai?����Wn
�q
2�f��l<�tF�j��)��h�������P�U�/�V�Su�Ćay�w��߭���3hy�Hkq��n'�v�q�"*��! ���u��4�\_����Wo3���D��ҏ�qj�^z�ρ��;&�ܺV?j�d�γ/o���w����NsQ�(�zBY�v��s�CTc����h����A����bI�-����~EwC�����W��
(��́7���QxF@��}�?���!�Ԁ�~�rC�[af��̕7,��n:�L���C#�k
�ͭ#��v;�� p�۞Y�)��]�1!�U��0َT<ǳ�)�N��Ox_bm蛶96&��[!����{�x) ��I5�(�� *&�Р��:�:��l+�ֈ)�v%b�?�ƺ6�/���H���t��Wb��|�&|�A4T�g��WnX��XNJ��Z!Bb�GL�c Tl�FV#�B���%�F�x��\s�i2��{�|Tc��p3��J=GW];+dY�u��`*u��荝����d٪>n�܅����z�7I���M5\�D"=�����V���EI���������/���[�my�ub�����*Ц�%�E~ɥ�E�7��rm�F�$�qv��w-=l{{�-n��B$����̃
��9#I�����|W�\������[/�2���}rC���܊���ĸ��%�w��r'��E:,�Ԩ���~�)kϺ4豌�_I-���3Z����y �h�i) K-#����<�y1%<0i������*c}����k���"j�k6��5g`~�lj���_��6�S��^���3��V	-be�X4�bG�󲲼�_蒀wh���P�j�K&*�a�