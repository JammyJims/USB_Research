XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����r?��K"�~[;�o5s�8��cv��'E"�_��7G~;��p#�rЍ�'�0�_ה��n���G��#�$�j���ٛ -�B������ܵS pP�.�%j�ue�x1�\A�ͻ��U�T:N`����S�Z&؍�c�PQ����/���K��3��P�� �I�a���[�V1�ğ����v����h�gˬ[�_N*�֗��q�:�Q�9_����p���X�[]�9�.q籢���&�S]G���q��_ZT�X5=�j`���ǉ8�Ԡ���[��5P��\ī�g���Gt�C���q��5�PVу�p" p���FW���;sF�#c;H�V/W����s�g+-!̀RP�<R8��_��X�ߴN,�^�^�d�B�GP�>$Jοr�;�""w�Y�ǭِ"e�~�{������y�1E��Id�ډ�0���j��%P�r;���xk�V;��S�O��aM��iY��8�W���*��|E`�ș�3I�$�9���4An[��I 1����hº��s�&�Z*��ﺺQ��?����\��ϡ�t��={����r�r�ƎM�t��b�:�5J���g�)����DS�b�,K�9U�y�w�l�ʒT)�P��g!��FS�����p�uŌ�f�%���lɸ��>�}�m��pYh�Zk�sg�e �W�q���4M��-�:�(���QC~B��5����ހV��,�˵Q��Q��n��;�}��:�������Vq����6�w�����5؃V[��XlxVHYEB    2ca6     970N �U���O��[IW�{M�ǰ$��nDY��DG�Xր�`�p?�]D7c���N�i,���$�_���������^/+L �!�:��n��Òx�
����%��_�Ww8���8��5{�;?E�ZLy���V�)|]n�v������ǵ��M��� ��@��܃�>��{���j��E�QS?ɖ�Y^?�:U?=1�*H��.�q?Ӳ;|�7���b�	�^;���/���]D��0n��S>��xѡ���ahH��S���n�i�ӊ[->
~8�do���'L�GP�j��zθ�R�������}�m�����nkϐ`\d��0 l�v���0���	j�c��ޒB�{Y���/w;z�+1��4Ųg8t���:�7#�\�Tw��R��-i ������̒�Y���z�:�=����{uЧ4�'��ϲ7��#!-�.X@y(ّ�u<�E��&���x\X�6�A�M����xzR�O�`��w�Hrфgf���8�kc�ln�3j~�}��58�՞2X�FBp���fq�NH�Ɗ<�^���Ep�gb��;C��49M����.�xD!��;ͰA�B�,&͝��m�H�r&A9	�3.f��9��i�J�C�"�@Nx����h[���!��[yjm�݅H�4��v���bQ^�%Q��E��1�/��#�d^N�����ok�����Y�m���	j��O5*�g�̊���Ú�-������X�P9���]���F'���ǡ�"���l߲T���Z�*��v�o���{R��RHw	�c�bkh�Cj���he:W$l��H�� 
xz"�����:\p{;�-�ϡ�|Z/Cg��mzǗ�H���ؽ�ϱH�p�,Skj�Z���3"@'����B<��lE��N�"<.�^���][f�RE��@wU]䕍�Ʀ`G�$ci}Ϙ'�]���T��u �o��>�?�PX��"
r0O8M̈́�,Lu�h��]��A�'�E���B2��+�v��VP�.#�z #,�)i��+�,�ݾ���&��׳��3~A�%�������?W�w���eg(�'�a}��z�T�w+Xj�'��A�����#U{�JD�J���U��y@b���Q]:�vbk�$W�g95����D�փ5f���%�qZ� ��u�F���tGl�)w�A�
\�:���3���|ޱw;�_DNw%}�.W�'`�@!�3���1W�S3���R!�;�Y	?�љ�Z�,U����r� �_��`�i-1�>wW
"�]�
��	��0I�uk-�r�z�j����T�{W+k�$> y6�Ƀe?`׈�q�/g��Y^��,��,���%_+%N�HN�:�թ"j����H(Y	Od���+}�X�3"�t�/�D;�I�w%t��T�qb0�r����\=kl�a�P��K~7�S�o��ڨ��f^l9�UP����dy�/�}�0Ee�=�T�e�/�05����'�W��lY�!���� �X�=�YTp5~ć5E����
~���Y�(K�o�.��,|�M>��r"�~1הT�x6s���Mc���S�����Z�X��ׇ�'aR������WFzS�Xz|/X���9��u����e"��D=_����D�}���ZԴ���~S<�6$:
���<�h��вM�h<H6'�;�I���Ϝ��
�3�h�^�nVsԺL���9sx��\��'9&�;�љWf���/ܗ��f��@0�G-J�H�g���#��BoMWK���LDvU�U%�hP�3sF����4��'+�<9��{����T0���)MW�-��u��N���C��8�-͍q��*��.��L�GPA'T���~���{�m�j�@	;�4eR�[��qX|��%����h�i��]U��������1��S�N���my��)P>�Ak���&�ڻ��U����^ŷ-���ؼ��Z�F_���W'R1�'$_��m[!(���[,�>�^\�����A�L*W��]�y��y����I���/�[b0XC����l&ﬔ�!1���ɝ\�O>Ќ�1�e��
)�iH�a�j��}����h?4�JUq{	@�ua�t����Ģ�$4�2VCO�8=ƌwpZ�Q�7��l4�]��!Af���g��Q�{��`'u�p��S��Q�
��/��d�����v5=�Ҥ��J��3W*�� ��Hԇ6�Fk�y���M7�p�6�����7�
�Z�ec��'�٥����IV*g�	��b;Bc��F}͛�*⹕!�G�"i�lLZ[��Ɍ��7�ྥ��K��S����C�9*T��~1�KM�_��'�i�H�c��+�e�$�m6j���.��Z��D.��Ha��P�7�'i1v��[z�E{y+�0_�����