XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����W3�"�	�E�A�����Jgϟ /�D�0��/j�ۘ��tBn��G��S�P���
��u:}9�GcV3��,�*2�	�-(aS�`��z����(�C��jn�/.b�F�Sћd�,�vVU�����Cͪ���n5P�$�=���G�%Ԥ�T�*+��9=J�}��O�uJN��>��T�	z��9���'i��I��i�jyT�<���Bը�yw�JϾ��t3����)�����4��#�e�*��J'�z���s�uc�>f���(�m���[��	O�'�sxx.�_8t ����O�� m���$hWkjD`��j7h���	���Ʀ��B��Jŋ�����z���>g:6�0ʉ(t1���!ݸ��	�U���mq��ѕOh(�}����:����������W��
!E���TXfv����b��<6�X�0T�3F�xln��,��� �B�z[�39I<���_��)�?Ϫ:\S�@�1�^�۰��3�%�JQ��V��"6���m���=�t��7Os~k4�F+{�v-�wqk�q�Ρ�w�� ,���^�e�fOBB8'�#�J]���謞�����a'��_A�'}�EB����2c���TJ��a�eP5�Xs�:Z�����[�mqy����#�U��8W�����_�s#� C���[�����ۚ�ܐ�<�^>@������Oj�ť/o��F@�u��/1T@3�
/i(#��
K�0��5���|��E��	�C"�XlxVHYEB    45af    1380���J����b�,QE1̠�Zd��+ oS��n���say:���������H=Q���lv�g�Y�QAc���X#78?<��<Y�xϮ��<Fs�S�$����I�zM�� �b�:�w�?~�6�J7�i�&"Eމ	�1����:S=�?~�?b#��]vR��
�R������kQ!�7�U���x�C�`��­���lD���#/
z��F���=|M�s����(2��(e��z�O8�|d�����[��.���U�<	h�j��-�ԙ�/�C6@̀U=�@�!2��g(!:�Ҳ�F�N;�~5�ae��sn�侇�����(/�iΚɟ���;O�I)�2ư�\�T�F����ViO��?~f
@�|%���7o㼠}G8$�몧cz���C״E|���9kR�F��t��u��$�d�������ޅ(��&��r���17�� �i�����(����UyK��Il��W�9׈(Nc���T����Ō�Ƴ��1���1����K��W�y��?��O_Uk��gz���t��E��VU������~U��#C��aAiՃ�'W�q��%x.�;���k�FvK���B�H�2�A��Ɯ�@�x���B�˭�构��P-s����!G�8��5�i�%��@����UH�Z����������[�m�)?�I�0`C�3�j��C�i����X�8Y�� ��mӊ��E�D��|r���D#D(:����Q��kخ:�j_��|�{R?����r<=K��/���^!�}�f+��
���{��l�K|<[�����%�0�Ѹϛ�Q*�m�V�����Y ���o������Z�^N2i7_��g�,���ýȷ<6ԟ�nk���gR�kZ�ii��zg�D]J<�Sz�t�ifp�{V\`W�E�� ��vo���u�kbOs`��W����3���O ���o�	�E��I�
^F�+�[hQ�E��荈���b7h����NY��)��B� b�.N��_�xZD�
�x�D4�3��|5$�"p��U�z�-���uI/h>�A���-d�],��(�-�!ٲ��?�-���U����`ݤ�����m�;�T/�=��"h�s�����O�T�9��4,�����5kZ�ꛍ+�2}Kʣ�@K�>��[_�G�^N���g�`���(,�N؎�](z̚�x���=:������"�GG+�.KM��4$U=�}Or^C˽�J_R�N�H�ˊ-���*�O�NMs�=ɯ>gԒ��ĆnA��s�/�#eb��9�pH���= �&X��6�����u�D��)FTQ�zDV��y쑺�4��S��R��e����;�������>Fig��*ôfP�3�,T�,uV�죢�-��1P��Ms�V�8�U����P.�F?�$����L-8��L�����g�畊D�{=�f]�?�9�1��|�%������6��o�b$Xm֬]�f�����P���|ޡ�A�)�c��5�|���3*���� �GW�ތ�԰��Y�������?�<�DJ{#vj.���b
�~���70�ҡ� M8C��&��,��	�qfu$�H@0X�pg�/��x�Gg�i���]��������>�v��nB������/z��;�F�@QgN#������Dܸ.�ʅ/�&)zA5[Q�4i�����n=ŏ�u��������|U�<���-v&��[�b��}��t Ƃ+�qSDɷ#���bw�o?�kB=~iD`۝�<r�:��It��������dN��.L�l�l�P�&��� �b�]��N��s<���_�����RM~�bS'��X���~����)'���:�ڳQ�g�H
����O�X�m���b7��g�8![��	�6o�A�2���-�)��!6���|�h��h[=)1�_?�Pq�����F��AMlCq~��<�%Op��r�T�-BL����?�}���t����3^�@F=�R���2�rnwúf��B�˝7m�^;�'*_0����Iތy!6��c�&�e�FZ@��[`)��?�C�_�J�08�+��OZ&-7���;
<�!�'�{����ƺQ�M�4�K@�(�P=�4��@�K["��WMl�~���8�#V���0<��q�&�?JU@��d�!���#���X�~���)��e�[��K��@m��:38��^;��x��Dd�'�$�:.�{t*\�GM	;K% �s�>1f5)뾏1��uI��H䗟�i:YZ}z!�WR��������k�9o��Ęq��
^�l�9�{���uKÔ�kZ����+4��Y�<;S�'N�#:ZX-�hW�ڄ�B��*lg9�н0�^���1)��+o����� �vE�d�K�c�~�=B�W~oA��P<Z6HR[�ם+�i��?=��i�U�`Y�t���Fʃ�{���߷��1�:I��甂��=xB��� ���Q+7��4��?�qj;]����p��������t������r�y�/���ꦭ����'��1���#�';����"X�4�Y�yn��+�����7�V2��S^=)T�udU �Ŗu�]R"���^�n�#���Dd��o����ʥ�����4]Ki���X������J�Q��¸kF� C���3#�?��-��_E�>ÊX��AH�}pu1r��t!�
o�ͨ4_������L�D�oقGM������V�Y�է�2�3!���l$����S�i��)$�qh.�0 ��43E-U,�G3c�F9��&T�a�-c	m5�PF~M�7����]����gl�jQsp�Õ�S�G���9ɐo���V�N��֌�����_6Ah��K24�>�JI���.�%>=Fr��UQS���2]8Q�2B�i?�O�vڂ�A<`l�:Z:%�a���]{�<]�z�������$�6J�x��M�wM�Sᶊ�v���﷿���]��8��_�/(�N�&/[Xj�?�XfƎ�o�[��l9\�qk�q5�(��ј��6��O!�0J�.a��m���#�?U�1]
��'�}�y1���e�I#���澳�Ui�m���!�k$�ޚ*�J�Yp[I���m�}��#��G��#=$��f�ʷ-G�wG�u�MG��T-EI�����1~�nX=!H�n�t9�/H� q�Ak2Ei�bN<��㑕ܣ[�{����	����v^�z
\�"xH�аab���/��Lo�C+#=ۊ����N�x&���jh��Ӂ>ԏDa�<�8�)"B��6\`�r��4M(�����N\�(MZ�f�&0gV������
G*���I�=cg7��y���;����9�f���N_��BL�tm�b�;%&��\7��}<k��s����A[��5D��O <#j&������ �[g��纆�B���E�X�;Z�DU���Ad.5��b�R�����Etk�B�d�}t��gUZ%k�gG*��|ü�6�]�D���[��=|a۞��4,���j��Nb��b���.r �;�
��T�}S_���(�T�K�9�(��okh��?Z v�F:�U'��N��F��X���F��ϫ�I�����Sq���Ke�K�pN�N�2�Y����I���$i��F�О��#	H'�T7o���-8<�+x,?��+��&��f����d���I�vǓ��:��x���	O]FA.zː��Z3cE�v���v�[�]k� ��q����`=��a����!�=�*�l��!��E
�H�4�Y,I���H��-����\����ɜɨ�/��X
[�QO�H�Q��v�jYo���0��rۜ67�V��t�P6�-��w��{�y��藬e�������+*�TMn�ဗa�֢ϐ��ޣ����C$f�k��@ԯT@;ǃSb�#Ҧi
8Ƭs�O�L���8\S5�4��tm�������u��UG֩tMJ��|�6�e�kxr7�P9����UW�� �U��8�, �ӊ�S��v7��
hDt�P�b�]��`�+<G�B��[�S�?�_(��^\�6P�C�*f���઼�*O:�Uӑ�ⵜbM؎��[y� 㻵1������\�ɏ3t-��h^���'���̼^��2��y��N<@W׷���q�3��]o��i��fbl/"�B�{�����)���װ�j���˄��v�(0���~��A�Wz�^q"�e�fB��|��>
��' �q��{�.c��O؈���k��M�d�u9���V����
�\A�zSV�b<�+,j��d,V&�`����}z�����eX"Z�A�c�����k�^�	��� ȉm�25_����中�Oa�ۓ0c���;ڕ��������0��J6��}{�u[�R�������J���ܱ/�m�$aa�˗?�]盿�Y �.|��ؤ��n����D��ω(���Ί��u�r$���
^��cVd��fv�-�ü?�fX�t���T�m��< �KT��������^�����=�elV"P_Pӽ��d�yH������8rL�u��_H����ҷz�C���ϛ��r�V��}j�� ;*<+Q�/�}�v��UV��DTQ���D���m��o/��:��LM 0vO\�~�]'���8'�_�A���Oc�qU�h�;�&�ET����c�2T�[��Ǳ�g1;�c��}F`���T,������x@��{䙒����� W�j�z��n����%�b���p՜�6��GU�I$�D�5B���m�g哑���8����!7g�49���,�Y��j�[�b��k�g���I$=���O層��˄]F�_���,���9�C1{�<����B&K��^���(�,�dfdX�\Z�x3�u������