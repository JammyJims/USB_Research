XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�tLuvluF̵��R�BZ�"ܲtJuTL�Q�s�?"�31r���8]�����~.�6G��͗�zv�(s:�{��S�m�KI���0�NaM&�Ξْ7�VcD	l��X�&x���7g�%�Y�2/��K�B��C���}^����!���Z����	�]�O�G�s��N�3:���ʼ��Y!!F#ˀ���_{�����T� xJCtM��lL'x�y����@I�Rl��F�7@�� e\���� 4y��U�s�j�&Z��w>�܇�!э�Bq3WfO�����{����[O/��=[��/���KhI|�uWb�w�2�	2� ��%��.�>���'�E�����A_oi��"���7�фл���/\��[fJ7vLg�ȵf�\|�!��������ؕK����<�z\D�r�;�f��Z��-*�jvA�I+Ca25bD-UEQ����� ��'��~2�u��n$H;{�jۥ���31��>EPE�f���
ܞ��,�LNl��_�U_v�� "�6Ҡ!�o�p�'5�����;y��7zRϣx/Vus`����(�W@G��yf���׽s��k�Fͥ�F��w��}]{�Jm��5 �#��S�*mji�(R~F�^%0�5�gWR}}��1�P�V�oܪǹuȬ��9y��3cU���t~��a��{&zo�U�=練�
<ѷd���čU�������6��=S>�ܯϒ(�9�"���"d�A�XlxVHYEB    191d     a00�3d=���^ax�4[�� a=���x����-�ƚ�Z�Q �`R�����VE�n�M�ά�� �,�L��O�oa
�ȞIb��\���C���5ԠW\EC�7C����]'��|1@�}��,�?�L�T�+�s����������}�"�Dy&��	���W+~Hf~4O�v,%��d&��N�S�vj�%��.L0�B�u�o�����5�$	�zԟ��%e���g[�P�8�#��Ht�&�
4)"�'~aM�S�GZ�2Vi�n��Z|����+V/ڝ���[�B���B'Cfn��A��w�+]����]{�����5$E$?#~���H��Xx��X��ac�;*�����}d�
���������xq��Z�J����F��s�0�D
��	�����2��X:/��ѫ�;���ɋ��^ˀ�/�X'<�r�񪐤�ۤD��Q�G��R�+�*� �5��WA<����ĸ*}��4\�4�����ȫX\,�
dP����@��c����rs$�Ib�I/+��p4��<�c��W�U����x��!��}���6��(�n2��n׿#��R��V�����29����{u��F��?%�*�/gM�l�Y���;k�#GC:���O��Ĭ`&��1O�����׻c�V���d��J?s�a�Q���a*�u�K��� ),�ln����$4	ԟ���d��&�Ȳ���Zbt�޽�X�q�6�bڴO���2*0�c��DMQ���n�b�Dw
C�Z���i��Z��?��o$�$K5�B�K~�(���Lܨ���)���
�z[0.x�U�Kc���E�^Z��3�"e�كS���w.��Ż���X��t؊��05�J��*���{t*n�5_���`؉������>��%*�d$�nb�[#g�k/Ѕ(�']�)bKzM=֩���i�!��G��rs�X����$�2K�k���x�;'2I�Fl2u(��v%C��R��㝥�� Ef�yx���D�Kѣ�3������|���!�B�g�\�����d?,j]Y�j?�y����`��xν��2=�Z�����QY�2�Y�܂��Z��QPfyZ�ON��Hd���#��w5��H���BW>W���6���1E�r�Z}G����dbB<���V�ѭ�t�DK�P˷PN�P1���@�M�l��U2�5�˵�ﭲ6�`������(F��u=����5�����0`�o�y�e��.��4T�}%$&[F,}�w���:�1K\�E�{yє���4Z�'�ca#e����n�O��J�{���G�v�T�S�>c+�w3!6I��T?f7����.��]����t�H�Bm\�R��?01绬��b�N3SP��o��eF%Én�g@h��:M4q4�X:&_Tj��~���d��í�`�s�)�Q��D��H�`�m�tv����*�vm���\��Lr�(,��C���*�U�����P)�kQ��B!�M�����wt�b0��g3�JuY���X�|�Qԙe&>�g�{֦�Ú_�հh�?��=�.���zOs1�S]��P��ag��e<j�i��Ȯ���u���� ��ԥZA���z,��$�U�t.T�#CE	������R�eB���������z� ��:tϗ���C�N�4m
u�˩bS��{H/N�C�Y!���~������)!o��P��	w�ưSפ�rྪ�=�-q�'�G87�d壾�V?�q��<,2�su)�u�E�̨'��o��n�34����fD	���F�͠��֮�N�(:;!9Nk�鳦��v����X"�xV[��O�O��jLo2D�Y�0����B��p���P�V���Yv���X�l^v������8����V�G2FN�:��z�,3�r��X�0`�;�N���?P��2n1o��G!C�$<8cCa،A��u�[`�����u6��W/�5�n��"%V�8KǶ���Gi�w��{�B�9Vv�s��:�1���gQ����e9J#�W+q���ZTڝ�H���!��_?]�7���6C�y�jB��C8���(�1g��-T�$U����S�jw#��9��j�T�Ƴ����{Ѳ��D4fSA�G4w����Ûq
��Gޞh8�jȲ{\T��>M9�t�|e��'�a�,�,��A�-�rt�j h+��4�0��*ba{�V�r$Ve�OΔ�YB?���b��I/C�m4�_��&�XA���:�yv�ϩ� �.�^y8���5Tϼ��z��W&��^0��x��*Bj"$�A|���Oȟ´K^H�.`��$ߩ�.T�T�UA�cE�j�#�Ģ�G�zLI�.귃���Z�r��(�����P<�:ښ��G�zt<F�`��b2�����a�,�8�{8\IҘk�F_�8��h`�xq��6 h&�t�$���^g�X����CM��Qsl�P�Q�Z����y�������`�'��J,�Y�%�! �u�#����\Qˠ�M��S۩���T�Z�A2Ljc-7m�