XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y�������Ԁ� J<טi�5�z�2�<���_�m���_�ǳ��A�5�Z�r�]�m\��@� ���kY���n�`���.����N���w������=�E��������fk[z;YcMռ��Ʈ��N�!��2�N���T��=ԟn���X���.7)|��$!+�"�;wi�+|��G�ƹ0�b]��I�]W��0�]VXU\_0o.]# �]mܥ�X~�����	3L"��	l�d_vh�#��a2�v�	��`���D��H��xs�ې�ٹ�0����3�����m���B#�俘����X��o�8�����Fw&��G1�O����UC1<ǚ�Ş��@1�v@���)�7�����,I%�Wy�a�o��܏~X؈�_X𓿑Յ�U!��a����[��1Ŧq�+���ҽ�Ɛ�9�	�z }�I�o���:F�c�g擇�$(���P�;��ů<���#\m�c3�W��&�X�Q��w��3�G��\n$Ƥ^u�DO��)Ν+���p�V���I�.90���GX`�w�����I�˿˺D���mϳ����n��=v��H���vpE��Kh˵�p/����h�F&+Y%2�uc$�kE��]r�	H��EU@ݕIޥ�_s3��1p"��'S��ZQ2%[z��b����������.*�To��4Tg7dL�C�W�p
6�!�3�9�_����%j�ۍ�������מ�`����P����o�1������Sf:�^1��)XlxVHYEB    fa00    7180�E�+iw�s���>�v�[f�nSy�q~�P�H�c�i���6>�@�����2�T��f�x�r C.8R䌲r![B:v�'\���#f���x��-3&���S{�lm1C������V�i�vq6�A_�[$|I"9+Q�M��2Z�#��Y�Y�-�8,���\��1O�}m�GR�z-���؇4��3�_+�Ch��2RC%9`-\��%e�*Pܾ�
�K��5�%�bB������Q��
<
��E�aWM`��vp�?���"��p���׎-�>ͿTn��u�C8�X+���:cq���u�3x}NX�/ć��.����Z�@���Y��q���<CXWÌ�(�QV���E}N=�p�l��ъU�SZ��7Eh���u�*���� ڢ��q�=䚁�ݍ<�r�1S<�o�?�5�9\���2�`���v����[�,/���R���@���֍T�7!.G�kQF�j͐2<�����Ǘ�|RK�r��v����j�5�$e�%��ӆ�=�>�hJ�|�~��V��{\����@q�c�l�2��V����R!��B>uc4R*��n��H�8�Ї��7��tFW�p����hG�H���+%=��]����˗����m�	g��"M���v�ﱇ*����6ȋ�9���w�����K�)忺���s6�ɓ"�tD���tD-Z1�+�x�gs�Sx�)��B�����29;��� �b�"�%l�ׁ+�2� ����J̚F b�VݫEj��1�� $S�o����=���g1�&rR�%�˳��:m�|�%C�T�"lu���!ޏ��3q"K(�,q���+q
�����޽��΃>���).9�hi$g�@��A��ۏ>��F�����fJE�)�c%��.-�� �5�: <����4��[C��.���Jfڐ�"9�s����X�$�y< YǪ^F��S���r^b��M��V�Q�b��J�a�y�ʳ�	�3�8Uܳ��ʤ��+|Z���X��ޞ���~���#'�8�݄�Rц�&Tr�|���ۺ����;�4�?*����iK�q���挰�j��1�;?��i��t��b�Cz2~��Q��9D5��:�%�¬�+@$�y�wQ�U�t�Y>�sf͹��(�
"z�>	r8Z��hq$��˗�s!��8���l���3vc��8�+�ڪ�˪��|-T9�Y��B>��Řk�N�yA.�%�j�e�A�,��u\ea��;*Kv�V�wph�V��{R��&� Q#�.e���R +X����y��(�yp�A�w�3�<x��U��OӲS�͙l�-'H[-�Ks�Va(��,�6�����<��w�a�NuN���� 6��a��}���B"�m��4�vß��Q*NLt�y��4 �����������-��8��C��^�LݮrML��ؿ�g�P�]���hʌBù|�j�K���`l���8��Uv�S�F�a�yJ/1�p�r���^߀y����Lmݜ,�E��%��З���9��Y#z�ϧة��F�ԋ< ��k3�%�e,�;g�}�E�9e�l�N�2r��X�`�>+�-�f� (U�K�G/�ʴm�n��9�O�DN<��f�xҳY�k4���5^��4��$O��J_���n�W�A��M'd�QX�Q[��J޶4r�/��ޡ@mbkq�],�z&*��.y��$��w�Ku�ߏ����Urt�G�T���y?>�����54ɟt1��:�= <�0�2�ɹ4�'�����G�P�.�9��BtM?Q��&�d��s|/ʶ-eX��E6�{�����fd��
~��
�_����2����ΓA/��K��a�z��X����$GMuP�&Tќ��
h~q�F���/[�;e~ ���|��·pa/��']O���19Ymp�B���F�� �m✯Ĭ)6�
�:�	�`"x�q",�6�J���$D�L�n��X��wВ�O�� hU�'��$�:n����DV�,ov6��3
U�����Lf
�����~G�?�zH��%͞e 2듀���x,�
�����[?��'�����+b���U����X8����fPax�T�>O8d�X��}֌1�b���k��� ��L-��z�`�v7��;1�,j^��<7g{t���}��jAޯ���e(: ?�A�K^�?h�ܲ~�de:��V==�M��[�4"���P���V'��)�O�H�u��;�O��c���o��L�1�����n���MI���\^�l3â饧}¡FM�)��:��� `8�g�z���$���wHSw������o	�]&,`�hˮ�-�	7�eZ�	�X�Z~��L�~ ���{���i(��4Y�����g����<�R�d(��f����z\.��� ��LcI�׀��(��dM�"���du�m��� �ڰ�.[���mk������B��*�b
��h|�?[9?�h�L)v
��Pv��Q�U��Bl�������9N=,g��`��7Q]g��a�wƄS�
-��w�PL����y˫;q�]�����l�T�~�~�x����
A#R�'!B\5�G}����f�/�����q� �y%�P�������B�/�u5�ˢ ����vi�OrP�k%Q�*�.�Y�'j˭ �#!Ԫ�J�����&�)n@r�JbLR��ڸ��-֌v�7�� ��p�.�Tc��[	ӓ��(a�g.�#oV�j��x��Ts�+ܕ�q]&��54��!
(h����%��.[e��]Ppt����B ꑗ���Ǟ����o�N�F�k9����s��7s5PW�V�����m%��T�7sf�Wϼ�?��҆p����/�D�#���EVR����=�3�Ύz�=-��U�&p6x�9~\T�ڪ��M�0�Lɛdh���+�
�Bȋ8������k*Ttǘ��4Kx�.�]�<�j��ܸ�[+L���MY�TƂ?���}. t�<�5��	|1���H��o�� ���2w@��dr�T��{��/�e6N,������扲gZb1���S�Aȵƈ��s�w��ܼx+/��q�(���-�Ei��G�-,����9�4k�r�n�g����m��)�\�/�0�x��rv?�Ĕ���{
�,�7ɜ���zy)��
��7~z�,@��𗅤��,��Í�)I[5�|Vk����g�C���(�	��`F�8��Ѹ�jJ��[�e��e�p�Ծ3=�'�=�Y<[3����=<�3R��׀�S��9��6��7iN6B
 �E�Y�꭫��&�t4҇�hG�����?Ȣ��!���D�-f�?fQs�'p�t�Ω��P�nǜR��s�V'5�ͭ����F+��>m�;CB��������>j�j�-���r��Aj��/n�ߍ��F�y���?��b���"D�n��յ^��>�U�\����da�7�C>Y-���z���ehٙ��FS�G��7z�)���������
���ǃs�	�
���7�a6�j��+]:s//pX�~x�a\~.�R!�οyYM���Z��usBm�ɢ��[}0$6m���ۼ��.X���M^@v�Τ�Ir�(�g��I��e7xU�oS�h�` ]�b�D�k����C]�̤�`�$l�Q]y��kn̈ �#���	���u�VY�E��U���B&�u�wxU�βa����l�Vؘ�\sD��^f�Ύ������ٻ?V��_h ��ἷ�X�y�j�Sx�}���˄�+���WV���2��5����$����X�:���D����]^�wޜ��I�b^Y�ލ]�H+��Z�$B���>�\��V�la���"�W_�1��`+����,�f~A!eXC�ůn���31|�%
M!�Gu+ʌ�Pt[[�]{�E�S�v)��cZC/ �w��[3}x���~��QB����tB�Ú`X3���b�O�ťn��I��MT_@��xfO�OÖ����� 9�X��@�$r��gu�cjG�K�c�;	#��v���d{��{�����X��w�C���V��B�F]h�r!i.�t	\xjh�R��<����Bz����\�6g`��ڐ���W1�z��`��:��ɸE�wd��~M�3�^ T5��x��&S�/yAw7�N�o
��J�?�^#�ٲ�~F�&.>���,}��\��4�IuW�zn��8���V��e�??�D��d��#L���t�5��K��$�b`$k��e �ʬզs�aox�B"vY���XL��ѩWɼ3"��^�%�/h,�Ml�6[�a1�s��M��o.U�������?_�Bp:h�����a��ܭ�4ɘCqA>b-�_���3=\A-��$���8��X^{�d1��o�7�Ga��q��*��P]at_�k�mL�EIg56gPX>l�\����W�vY��J��N��1�x�Q���6h\�0����E@b���	`�T<j���v�O�F�S��u�M��0���7�
Hm�P�ۂu4��,�.��.���t��y���<���X�!l+�55���[
J.���Ye�ߡmez�8��d�<}$����k��݆wf*yus&�=�� �������=aeIȟJ��{!��n!�8#`�?]')u�;��ܿ�yX���TC+�Y���2r<f�߾�8�1�|5m������}�ť���Q��t���Ԗ����g�b��]� s"�mK�4����8~N*�!1dR�2V"���g�<:�
^y���r���G�I���ɔ��0�@����䱉hB�*`��ܣ�L�yҞ�5�su�s��qw�q!Ff�T_[&�@����K9
t�#G�ɲ� U����B�i����,5�ܗ�?O�lN������a�2�B�/��˶Y���H\�,�$��Ǔ*Gs�1�� -�Eu��B���A�
��f�p,�:�[��r������H��#8]��~��2����ފ�}����^�ɚ����LR����r����R�q0 �Ï��k���Z�}���/�~j��ܚ{����<�6ķ�\�)�ZF�͡h����ݖ�Z�Ϲ�amQ�p�{�+�-�V�C��$+�':M:<����0U1�%P�
�;t-���#T��R3!$�����Pl�-��7ȬG��N?�A�5[k�n������$ϭ|�b�b�W�u��X��E�BV�z.�KȜ��թ�"`O��P��T�b�w�I�dVm �Ja5/L�����Α�ߙ �O�����JT����ks�?�U�P�T�8'�e�n��0��p�٧R2YY���2��Ő�6C�G��ٕ_Љ�8|{p��I����k���.7�o���d�2��Z��;~�Q��:��bJd�SFT�������nr�jo�ى�$���-����+f�!����ԥ2����N��A��1�'���g?|�l#:hF����Vwh314Be#"� ؓi�F���A����g/t�VjZ��q�c����C
_�|#-�~Hlz$\��DQ�9�d�Mj0�N���c�ɏ:�V4|b�K��o��c��4�+�O�B��;�3��H��Q���?����PeF��x�ƒUuko+�*��%�TѸ1Ѕޟ�r�r�G:��pӒ��$�|�޿f�yQ
"�������ؠK3��kN��X_U�>���]+�3H�z(�����tє��F���B�B�~
�VE;���O�??o�����J�Ξ		@�O�c�J�͞bY�:؞�i�l�Pml�i_�%X�kqJ��pC��G����t��Q�CH�HMp7�A��r��N"\�Z�㲷����f
�#��F�^��RD���C#�D���k�e��b�F���&�젏���<��\��c^�j_N����
�=ű�����~��vJ7[l�<q�N{�4�T���d<�7��)L��7�C.�;5��"9J�����,F�PN0�s���U`=P�Ҏ�nt���U��ð����	����IR?���,������F6z���MR�d;��cҦ�yZ}����|���W�)��c��Vva��@����׺f�
��i�uT[0K��s�Wv.��q�h�Ӂ���3~y#�[�׭�7@�}�����fej6���қ*����`���
�`'2���5����a-��Pg֠1�ad]�:(OF���.\B[�Ӓ���v�G�^��??����,�ƈ�c\��s����C�ҋ���W�8�&�=G2�qܐ092	��A��}������Y�]�d~��@0F�`S�|�b�y���db�D,i�;J5e�%I._w)So��Kޭ��<�õ"�~����xw*L�?�q�������pjM�����w}��1�:��AXO$q˅�.�r?1��Q�2E���<�.]�H�x��9)&���u�zLo��!y6���I��L�
����mo��n%7�/��K�1��,A!N�oB~�N�K��������D�`A�З��u�ģk �>}	6�n.������j�@V�ݱ����m�'F"d�^~��p�Kv_#0u�7��3+s�=J����l����"0i;d�yB�CV*;6�y��~�e��k�j��f
�����d����� a��g�B?,V�)���/���9��^��=o\�A�l�!G�n�C������a�ؽ��� ���d���R���:	�	s�{���Bc��%"�m�Ӯ��-���r�4`����F����ů�X�����#��Ͼu������Ҍh-���?��z�0����f�|�w�z{B�gFxf.V��(�`5�L�F��+P��~	�x?Q�!�C@����	���/qd�S���gw��Cنт�dA4,b�NqO�U�Q%�8�N٦�F���yhE���ã/�t���'��S*dKF�J�!w�YF<53�y#�~��?�7~��d� ��j�%�]�Q�C��YNo�R���ɇ�[���\�!���_ٜ/ >�`��d�!I�sw�I��;b_щ)�++�������:Q�C�t������Y��r5�_J3֤U].A��
��cQ�X{�T�'�m��5��?w9�Ď@v0ؼ�<n�F���Ld�����V��~������!0��Coν����U�L�ϓR�M�h�Q��%�xʜ�RK�<�5��aD�#��^�� ��J)/&Y�IjUū*�^V�Xd�-�+�C���� ���7���>A=���
�G�|E�v`��Jt��u���?���Yd�rM����������s�O�ȼB�FPL"�B󝌄�Qg��LP�Mb���Wz�qۜ5�6I�'�|e��_�ڟ�a������b�,cv��\hR;����H	��V���������\#�F��7;��SXi��H��CL�Ќ���]Hzc��˲�!�qrԄ��d�j��� p߾�� ��O�0��R�CH_@R���~|筃z&�p�?���L�����+㉳�X;V�k���@�H�'�>P �]�B������]qkĔ�L����D��0B�Q���,*�����ɨ�@��Gy0�CK߇d�#Mo�`&��I6���5��?^����CcL{k�)~��@��יwK�m���l5J ��Ë<uMp�(���#!z6nYA5�e`9*\��O��q���U��vb�X+_w�9�I�#I��Ay�g�t(cD5��RmM���qꩌ�%��\���7�Z� �J��Bôqv|�'����V������d�M7��U��޾4-{��-U�f�_������u_����R��R) ����MlT ��c��G��+��T����x��c9���]`
ES ��MB��,K��*��g�S�}�����������3�-s�ng:~��Zܩ�� l�I��!%#��W�����b4<< ��[���L��%[�$���hy�_a<D�7�L�h�1���j����7_��]<�?����f�>x���:)������c���	�䁲&1�]�4Er�8=�H>�(��r��� S��:Q�s_���H'�ߞe�-�]4{ت�Jݗ��v���Q9i��TX�k�'/R�vYfܵ.���x'S�l�����&�c�]w��r��qR��X����*�����3TB��;I�x߇3���	�d2�B�R��滧��U���8�?��(�����|C�Ab������o
x�n�mj�O
��������Hhm�?Y�%�]��!J?RH`M���3��Q��j;�����!��v��)����b�k@RnX^C���ER�)o\��<OG���|g��Qj�\�{�dh��!iՒfz P��w���D���"��'�{ub�,���s�$��_�P%���v5�TW��4K�WUW�3Z`Ԁ8���f�X��Ic���	�G1%�=$4$V�Şh�����g?�]~��h��#;Y0��|�/#��8�@R��@��S���=P��wU���ϿXٱv"��������(	%E���!�>4��%@iB����o#܏뮠F3��#��[U����VY��cjxwW�D0��$��ij��n�&QP�ѴH�*��.��s��SP�]���^�C��p��{�o�0�����qF�(�M��O%�0x;X����LyXޞs����$��㸵�R��j��y�ͤ6l����&E`#��yM$�̏�zD�0H� j���7���
�k'*�o�Џ�3,�=��.ڀ��
���`�#Oq��²��1�n���#;pa|g:Q�n�L
�MT!o�N�Y��i�w���~1��ܼ_]��_c�J�T� !���"��o[�'^ѿ<Nvz�� ��-ʅ�����Ls|��W�39�Tc��4QȤ=E��$Z��}'�ɷ,�:�Ws�u�]�v����LIpt�}��T�A��/�zj����FU��I�����J݁�/:�Q�6׽u�p�� hU��4I����<KLP]���VZ	Ç�i�-|�AQ<{�n=��v�ד���6~8u#m�k38%�o!�t}rG�>�4B1���3��0@��4�_�KDY�9R>٧YC!3����.�����Y�3��.�=Ǜ�b�sPr��3�Y��%[�X����[�}iqK���^����&t^�U�5����w��ՙ���2%�Q�$+n�)�i�+7��6��F��d,0�j���j���3IT��@��:+�a�(0�t̘�ώ��f��ώ�[DBA�R̍�H�� ˛�q
4��2�ۧٯ/�>��rw}��r+q����vh9�<(��H�B{&�>6�+%���\�����D�Y��<Q~��t�x��M����㱛@�pJ/�`�?3�@Gǌv�GNL���!J�'����<s�r�!�H�X;1���~0�����u��2Ͷ���H�9��"�Q4_��C�iH����2͓.�<���?�c߻�e 57��d�Z�^P%�e�14�З�K��g�/��-�ڑg�-v�QЬ�Z��%~a�{�NC�u�'�Tf[���}3������,�Q�D�Vx
�l
)8���M�Bz�5܊�u9o�Ж��"��Y9D�E7ȸ��i��~��rٽ�O؃�����'����q���'4��K��=v�� 3V�!�|B��w\'���i��['�7�_RX�(OYK����������|�"p��\����J�r!�#��(Ø�	Ő�>��N`u��;?&�eNuC����oh���f��ע;p�*�`ׇ��5�G�ꬼ��z����9�<e�\�7��z������;����o ���lf�JO
+���=:��'B� ��^R�&lې��Ҏ��=�y;{%��M�웯aRaT���>�#1�C����q��	���9�7������p]5��%CG��/�[�K���H1˟j"K��>&;�2�����|;*-sΨc_�YNai>���`�V;�,`-�5KC�I�'�Pi�@�L��d�AU�Y�G�?�}��+�2h��'�f�F��3����0�&��O,f�0�j$6�!3,%�W�����4�OP��m��ߤ�h��qb�E��>�:���=���;!�����6?(�U�:x��Sm�xZ&��E������³���(���eY�	i��[�3k�֦(ε��{�_>L�˄�I|.pҕ��b�s�>\��f7)�� �{:	��r�tE,�%m*�v��A�!+��bs�R��7�y���}"#b��*Ӊ�f���׸�>�t�@3.<!�K����{�T�E��5
��������vV��Tu�Fbl�8��9��.���PR�<���p��@ZU�S0��'�4
���'KjC&I�<	��᯾{�,��V9�Ĝ����(5Я�!�L�q��=t�h��y��?�v�nVHU3H˓�r��� �Ȁ�4j5wV)B�]�l��\<e���9�뀏�0����Qu����Q>X�7�i��퀉�����ލ�\�@~4�ݶ�½_Y�|���fv�x��FKOV)C��GSw$e1�����#�"����3~Vvg�c#��C���^��v�!m| �[�6�($H�	�u����7D���Z6����,� ��=���iB�#S>̎�[f5�%Ԓ�����i�z��U��))�j�J���t�%S�G�+:Xo�jL��S�,)����a�^Ef��j�u��G6���b��M�uU��S�#���B�aG�v0��߉ϸ�䴐���n�`܉@ρ�j�K��n1� 9ͥӾ2.���*�'%�X�:�-"n'i�!�񒂛qMhGF�hf�衛�1�L0M�t)�m���x�)�SpI+m܍Z�E��t�c�kvN)�1)�_~j͸�SyoK����:�rp�5��`��/��7U�,3;X+�+�\eO�G0���V��izAp�*C��2����ю;���*��m�Z�Ϩ��y�5�(�9�,�[���Mx�����4�I_�PԔ�=��W�Þj���'>�ʶ��B��C[^Sf�ҋBg~��,��@=P�����9F�'�v�N^���B�9;�A�e���/�@�/NE<Bs��8d�!�Cd2��O O�$��Cߘ<�-���۫{�#��yԗ�~q9�~R%�>�	΋9v�� ���L콀����I�n�g�M�bm!��S ��{SW��*���M2���<X��$�2���?���N���p�%�#�'5�ÓI�[z��l�����R�X��>7�Jں�z� v6惚f+9���(P_w�~�0`�������U���P����y�I��y��&h�R�(A�Z�Κг��v�ߪ`�̟K���@�Ƣ�@t��2��l��V�3�}Sy�)T%>�nC
M��#r��Ky�ؽ�\��y�Y47}���cS����D�]����݄��|Y5g���:Z�8	�;]�\Ң�@�ڴ��y�,�e��?���V*���T��A��8��e�2������i�;�m�Y[@���(�0�=1H�N�T�
�vt�=���V(FYT@�	`�#A�j�� �빙�xo��%g�(<� S�k�C'Y0<��z隄T�u�ά7P����S�1m��������qæh<�k�����/���	Y,�S��~���ǔN�ٳ��Z�v�*H���#2-���5�� S�z��0M�N߈���Q5rQ�z�)�#�ݿx�+zd��~` ������H�4�K��)���Q��'9��C��J��1CĊ�w#���L����#��/�.���Z8��+Ü;�.:�_�����o����c�8?��㮌�>o/���<�B��|�����ť-){�q��D*�:�e�i��SQ��|"�ЅHH�4
�i��>�]:-C��O��k�D`E�{�r��ئ8�V&�t�͈t�:�r�9���X�^�#�e��xP��Ĭ���0=�TS3�������6l\�+��S��ʢu��>��>#G���l
�}Z��_5��R�_k�*�sn��k���̓*��G@���E1_��bK7[;CY����艥-Ջ�3W-�ׂF랫��-\��\���ٟ�NJ���GI�^řSY�:�5�űJ7�^���a@����Ʊsf�_�I�36����>KGQ�!吝x���N�{9צ�-�B�~�e��N�L�s�"�}怈���r�pio.��@EP�9��:�B�⪧��l������aO�����8-H������c��\< t|�a����Cɞ��q�6,ՙbP�[g_-�Jh�K���CП��KK�0� ��L�1�8�;`Ќ���.�c6pu��ő@�X�Ͱ�j��Ԉ�|�J}~K�a��R�'�=#( �`�,�6/�W~��	3�v�:<��q��t�SeЗ���>�
7�N/#r�\�����˘̚+@���·0@�z��ŗ���a5�ۋ��~M���gbc��y��;
p��+J�Q�5����\��,,9���$��Eb�K"�0�`s���g�\���/����xd�xSv#��@,_�;ܶ��c�F`جՍ�CͩI�|c(��RH��P[��	��u�D��EJ�����*	'zT��h�x5^���~���3B����0�S��p.�b��7y��F�䛃ے��mlO\��+��uC*dXx�~����2�!�gv��`��T��Gނ�{Oz/7^�	��� �0��*�Ե�>�Ѕ
u��1��nߥU��w*2����8��`ӑRuHcj8�E��4�p��w�����(��C��>]�ꍇ5��#|�ҫ���Z][Bͩ�N<c�Z�ˇ0�K��r��J ���'y�����+���{<R�Q�J7���=-��vUqt&��+&4�E���WF������ �.%0'_MT���[@k����������=��~��H��ք�W������#>X��G�xp�Jfs��n>C����յ�W�"����;s�M� �gSe\��1�%*s<�!����� 6�_���,��f���6n���@�sW��`urqciF�W�'/��j�Keb֒�?�_��^C-I�m\���_��F=�Qf���_g�&1���X	�I�j�E悟T�5���p"'V�湞
b ;"(z['�I��4�!�=_��G�]Se ��FK�Y�hG�{P�r3���yXPܒ�H��,POxTd���İ�h�>_�<�g]�/.a��5�MV���Ly1����n�k�-V�����Ս��-5vBg�/&��l`
:�QA�~���4L��'G��$�]�?���ƟK0��IR�3�g�..���o9�G~��$??c"ܐQ���+�!ݾ�9b$������aa�p� /���a�;��"���jͩ0h�6�À���F/d@�������p/�ۥ���R&���Hqw�{��U��P6Ba6|��R�c��,9V�5�[�����I�~BI�U6e2��!sk��D��|�Lϲ*ś�3?� ��Km��j�C�>�Q����4�u�Y��u��	���B������e��vZ�z���FƧ�})z|�*�9J|!�7Q��ݒ��(���$�#r8mXūcߎ�����1d��wѾ����U3�iR��z��v���)��F;���%����J]?4a�fD�w l����}�%u���5)���j�ɧ�����Qo��"��oK l���eF�٥�:H�?3޸�)���1�|� �-D�#�\c��>i�т9d�5/W<f�9��.gg	��r-����.��>z�0��4�顴:�T4綎B�bM�r �(�#hӾq<lb���^��$9��N�j� ���\�^FVO����wv����%�#s�d���b�����4Ͼ�r�G�T	q33�.���ޗ�jK+'�k�m��N��[bi&�Y������ѡw�-���꧕���� ��`U�O�����4��\f"ZY���,��čgt���3&z�������B]�
�}���(36���#�#�h��%L��}��9D���Ԡ�>�P}p����3����J�s���X���E��%'�W�ݪ؊p)tFp'*G�� W�b!u�ij��~d���U�ĥ�]>rL�$�n,�C����rRY�)8Lz��x �<��e�Eg0ii�e�SU���������W�<����P��m��W�ѯ@����bl�Ѓ��[�8�#���.OC���(ݥ�9��y@��T������$��Ԡ���x!��m�`��$�k�a��kF�N��&>�j
VD��L�e[��XE���"����󬚦�5�i3⦛c��s, �5&)�a"7D�"������"~˘��y���\�u��Åg�r}v���ҕ3cW?��fW�QY�o������>�gU@��)}4�?*JE��J9��:'*���Y���ͺ�Do�����!����TB��%e���y˞�{n�qUҞ�ScƓ�a)9{^�ھB:�ծ\��3XQ� @�$��H�t!1���Ãg�4xh�[�����y��C�Dy˱mű�" (�H�Xi4>��I�h��g ��7
�R������a,�������,v �����?0U� ��2(8�儺�� �l�D�e\oCA#���5�"��"��^��(�t���
��6�t��";�v���
�/����3B*���������ES��5X��DPÕ%A��*�Q���Q��\���i�?�5�t� ����-����P����c�jo�-�"����m��[}.��)�t���ORp,̬a��2Ď��\:v��-���/�oAu~D3��G}-��ǖ�$p������#tY^�|�_M�����G��\���{0h���&,�Z��И�<��Q�9���N��j��#2��i߹�$��0Hl��b!�=�[��LI�4%��xj���(��x
���d�������PhrNg�߱�r�s>���\\��
>�C�Y�'�;x:!}{>�.�i�������&|��ƈ����??҆J���_�ka�ޭ{�y5CS�]A��l޶*u���Ng��i^�������pHn�r����ш�,$$v�8$G�> 0߫�Y�6^�o�[Z���KBO�Ԃ��p�%��,�(1����w��v8]���)�{���o��bf(���Lx
�U����@�eq!�m��ڙ�&&�3�����Hխ¬���޷I��	���ԁ}e_����B�g�q#x�g8�=Ѵ��;V�P��0��%�<��T%lq����<��Iǐ�FCD{� W1q���ن���S.O��v]I	���é)ܵ[ ɻ��H�/�us3��H��p�Eڦ�&��#�CZ��˓�R2u ��bi_I2�
�4-�F?D�5h��-���T6b#BZ��;p�T���̆�o92qjp7h_b��}�E���?.��E�儌���ä��Q`�d�̹3vT�T�����r`�K?�,hTT:�5H>`O�������34I�3Sr*K8]�mo"�O�+��h�,��?�U���!o��IP�����-�ꧫ�A���L,ah,�/�e�\Q%8G��� �?	GW�T��:�#zܭ��Xlb��G�c*����'`�th��81`3ᑽ-
)	��`��p�<���;����\����`Kr"
$�8|��&��@��	E;�~���W�4.kB�O�%�E�z}���#1Tw�)�q�_�i#»�Ĭ&+\��"+��^s�S���v�0_oq�1��^��;��Z$�C׈�����Q�d��%U�\��Tq�N��W��7�C���t��m�A:+�P�� ���c�k�Y"���7�]�Ps.2�D��r�An���'f�U�WÍ�'���]�>�"T����_м${;���v�h<����� ��pՠHM�)o��OcIA��Jj�%0�(������Y3�/�AJ9�[��>�q`�=z!=��t�����br�7^�����.����-�N70HW�R�ʰ��$b\6�-� �пgX#�-�4�ǎ�U���R���*&0ɠ�	2��Y�Qtt�!V^�?ת�(f������ce�L���A?�<�W�aw��K$9C�9�s�D
�x,A~�Dr�|�����=���?ɠz�%X+ұ��u��~���2)�8��+��X�g�tԬ�u���Z��[E��p��i����L��J=����]�*��jZ�V;��h�HH�_��wg�8��!ް���@��?����G13(�ǒ���8+��4����u�9i�`[�vu~�y@S�Q�X��qS?�R��Nuo��l�S�mZm�Q��<�*e�v4t�'��wSɌFx����J�����U��6�]�xDh	J1��É�Hr�/R��~���z��B�<����y�ڽu؁��A"�l�o�z_�l&���F�ݳ{Ǵs@��M��Yg7ڟ�dd�����؄�o2%��q:9�ՠ��E[���Ԯ�ɺ��\X�0�{��DUݰ��(�c��rޮSn;�.�g$��s*�<P�"
Z�v��c�E<h|h���B��y���E��}F=�����Z���a(�g GZ_�EDJжqݓ�r-�'N�Y7Z��n�}���CG�X����� ��%�x��`���i
q8K};3�(�<���
�
�k=l%V�ހ��I�۝^��]Wl����jT���Mi���Wf�܍e�v�dߺW+%�4��E� >�zD�hDo���J��av�}�%���GX�~c);h�P
�CF���j9|y<z����Ǚ�nj�;e�2����	P��\�=�rF��-��^�^zHr�� ��^��[���H�"Xܞ��h���Vc��N#A@5 m��� *�*߃��qc$���}�	������4�8�8(�:Ojg��5o��w�䣋^���˘
��~tɼ=�鞞�L�	�7��t���
j���+��oy�Q���=�\b�R�q�Y��j(���I�;ҝ��$y�/�O�1�ʕZ�k9<��ֺ�;������
\��kS��!�[�ǣs�RN��T�UI�&�bom�sJ7�Y�@�G^ꘚT+a7C�c[�d~N?�ׄg���?��c�� p:i)ٻ ��V�<����=ɦ��m�T1Ec-H�\5:�A��/p��|8�Qy]���P;��*���Ƅ35����T]��) )Bs$�
�9mwR��-6���t������r�z�R�6t윓�e%�5$���_>:��{��.+zJ�~���|�8��0Oo~jb��,�9=<��SD ��Z�s�
��R��~6�[w�R�\e84�c�Б�UZ��X�?�ֆ[�Lެ�\*�@���)M�T�,>����%�,���_~u�Ypc�3���*]F2�a�}��Q��>��i�)�1���³@�^�4J-�z�N:ө��Ѵ%�'A����
�~�G���V���uҰ=�u����+hsY��v����w���������R��BS�yW� �����߼⦅<��&+���y��i8�`!D��2��c�j��
G?�v<;���~�^QV����ūD�7�2&�$�W�ʘلȴ�1�H���*��b�'���<���^�����Yj�0�͸9E�8b�\!��{jI:ZM��AT�O�v��ʐ��,罒�kn�e��4�Un�~7�,K�wq�_�Y�衕e�?UiZ�B�N�ka7��)�.7���L=�ٹ�ѷ1�˳*� oi,��'�8��|Z��T���"�P�s̎�	u��
���^�	��`"9V ����Ў�?xD�#�ґu�xU���M��z�]�jAJ2sz�1X�����w[����s���3�	'C�L���)M�{7EpU�n�XѲK�St
	���~����c��n=R���T��F�U��(��#dγ;n���p��]��*.]e$o�[vP���&�1�r�7O'�zj|4|z�>�I�im�������o��l	A����7\�d�\���׮�Q�f���s5fs�(G����)Egc�9Rզ�?��>�� RW��oп� B~/��OM�g�����3��jQjg��.KpÆ�]DJf�Q�K ��px%!�����p!.�V�`�(��ݥݼ��!5�R��応����+\i�Ԍs>�
���J�W�4�}9��녘+Tϩ�O�xTӅ yAGN{�7���xh{o�<�
�o�L���:V�Ͱ���%#d� tV͒�ݘ��f�O�B����z�q�b!ʚ�W�d�Uӝ�G�E��>�x���0Bz�b�"���-B2�ni����~���)����x�q���{��$å�ۋ,����$����4m�F���f��8��Ѕ��PژF�5 �KFVD;��/�����2��V��"}X �duf�ˌU�U�c������7�s�F�S]��y����C������R���/m�4��!�m��Ӝ��en�tCp��\��2����Ks��a i=~�H2{$��z�2�kmH�%6������rTR&i���Jpi���um�y�����Z�M�GQEG������F���P��'��S�mkH2A��7f0�ј+-fd�rD���0�w@���\ ��I���$j\�|~�X�
�ϵ[u0C��r�_�i;����.�,WE�%�&��Cк2��xˍȲ�&m˱{�%0��)v$�
�������<M����1��%X�!~�u��;����� ����h��HXu_kn�Ă��~���1t��'tCɜ֌a�o����bO��{��.Q���u��W͖ip��,��w=c�JJS̙�L��{9����0e^����e]�&Z�A�׊D)|5������rj���؊����i���i��6�=���@W�֫8@�,et	����O��(#�L��>����>h-z�Hƕ(�/-B��	O:���)̕��F���5��a��=�t�!Ͼ�|�fi�m��c��8��a�h�j��!g���m ��9-��T����E`�1+,{q?w�v��5��A��g��S�Ta��+���X���m��a��ȏ��8瑣��G3�w�a���F)Υ�n�ĳw��eGs.ǩW�:�_s���S�:���"��L����ft��z�`L�"X�!Yf:M�M6��G�r��5co�2\��OB��f�n�{�ȝ�Y�Şч��E=Y��aY%p0���gb�U eR	Ŋ��4y��nK�����2W\�Te
U0���(ΩF�8�iu��ac�H-�r��_������T�&φP1?z2�R��i������<�0��z���r�V9��{g;b/ @��w�ym���"�#(
�p�_3v���C�A��kj��بa������� mbk,�������r{-琴�i���I3YY7�\������I�c�xh�ͪ��U+zM�|��Q/Guejl��ܨ����u�I����`F�\���d��s(�_�H)Ma������F�P��<�HS/j|�&� +Wr	�g��������	�sڛ�Ðm�+���5}ld�L�2��ì���f�X�� ���˓����Q$-E��k<�S����o}yۢE��}h>m	��W) �����!_"(�-��$�p�h.,��6��La��"�1�~,1��G����iW`+��D�)��W��Qt�m��o���������X\�~�-a�q��o�U��sq}�rg��f�[���<��r�IS�r�jD��B��`����>{]��N�E�\�9W����;��3[���W�U��=�p�{�����,��2A�'ж� 8^Kmtuλ��d�`m�8��B��f/&0���X?0g*�ru����Y"\�>���c1���G�aD�l��1����P��f�H<#��%���`�NX�[���i���pi'S/[��'Q[s#�^jWs�L����_x��L�?��v�^�k��f������~��P~d�c����M�A��2�Rv#�M��f��`&7Ѳ~���8����Y��.�E�� ~2�(-`Ѹj8�˛Ko�K�o��9{e�Y��B�{��G�+Y��1B��+\x2�[�i(�a�j9�S@�n� ��Qm�th��	�?ՄB!UE'C:��`�)I�>pǾ�T�^�d���#�Z��xD�ey�%�r.�#��P��l��+�H�׫��(lko�4�W��g|�V��w���V�������6��{�>@�_<�S#Rȿ?ƒ�FiHx��AJ--�5x�jU��R�%1��v�6%�7oM�մ5}��~���aOO_���͊,�ߘ�=��Һ�8\�.-=� ���u�ޘO�7�����o�5�u��hU� ȳ�&�t/�_�|+�&m?'�ɍ�ly���{6�	�de��EM����?��)��{tb�ϝĞ
66�?SG����3�.d��9�扟ЃMcOVݭ���#~�����wyV�xʳl9���t��~}�Wq� a%�x#5y��9��//-�LBXy>z����k�E����2�o���1r��@A9�6oI�/ٮ
��7�ڿ
	lg�(q�������
�QC� ջ�"�V)�c(]Z�m+�Ӏ��x��o��OJ�y��j�6������]����W�*m���}��ٽ&��}zp^>H����9�c
�Hn3ч毰Hc�o������܁8e��O�!���}&y}K�T�[���)��{�n��0ݣT�GR!1�`9�Mt&��R�[���vB7Ѳ2C���rd��o �)S3��Vm��W߲�9�x�����8��j�,Qq�?���o�9�ǂ���~��ҟʡ�)�r	3���U<�ꀼuP�����J���I9��T��"��y7�|�r�W�:,���[���5M4C��%��>a��;�c�T�3��{����I��*��%��'��&���q�E�B��rw|�+ݎ������zW\��0���_�!Imvv�K��&2�{<��'ɠӝ��*�C'U]�;�HX �\ ?*#�r�Ri+��*J1yf�u�c�A&=
�s�?��"},� �6���9iX졔�~s�<�&j����m��EU.�}���ގj��ĕ�E�o�ƭN����y$��kl����6��[v�]����Om--�='�[i���l����\ɽa�}cX��O�K�}B5�_���df>j�f�@������߯�B)�r^�*���8����/.(�dʤU����e��2���z8*Ku_����=C��Z����!S0�T����,��m��
X��'���B�	׺N�Q?n��8�ڷ�=�8yW��x[Nbp�j��Ʊ��߫3�kY�U�7�I���d\K{��Z��Zo5�/]���d����q�z��80��;��� ����g)�'����?�ĸ"Ug$vG��81,Oim���ҁ?|g��T��5���u�J/���2����~��&+�n�mɯ)f�q�h܄��o���1�6+Դw{��� ����䌇xG'&[���p��^/�n�~�s������{ �(�b1���	Jl��:+��o��[�5�[U�s��Bw:�^X��~��Q@ �ەa �z���_�h":�XPA����]�3���(�S��]�s�8Br�0<f�1��8��ɦ�7G#�$�&I���.��Z����ObP�r (,LP��#{W.���е�p,n'*(&SM��
Է�Ė24�V�'K��O�5�aF�&ҏ�}W2x�w}<��PD=�����{u4H:��chg�~۶|ɝr*�R�('�)�' R_�ԛ��+�~V��R�t��t@ބ4��G]D�b�~�V�_����ɜY��W���,� AG�F&�N��R:��[Kg������)��y�q�/�s�pf�4�(�Ư���Pw�K`�.Z�����Yx�d�9c�z����}��5��)N�H=fX�$�'���p{"�Qz�u�5߆wλE��S=p��s��_����	�/���3\ A�>�fH�.S#�A�3{w�B�4(Q���j�L�dT�����D�����֖)g�`�AA�7U��`cj7W��V��`+���M��{�
Cw㭻�W��79?�^Uc?�F��M�p�P��\X�pj������"���^d�r|a�E[{t���P��Y�5�JZ��6;)�L�t��噂P������W>��C�/E�D�I?)��u'����s9hծ�����T�1	�|#@��[_YF�+�����q �12p�UN��\ $_�R-�MX|r%`f���Bf��ɺinf`��B4,�0�F�N.�r�U�E�B��w���S�K���Ej�$������.�(�OaX�:���%h�a�k���<]D��4�e��w�<�2�=�h`�%�z�Z�1��||�F�+ԟn*9Х�����?��3f�0R�>j�c�D�B	�4MP��;�4���Lk��6P
*��vV����lN͓�L ����S�&m��
��m7#��bZ֯8�^��93v��m\n "�
¯�QG�����E:h%�7/x"���>����q|�<[��6��R�Vs��HB���� nIv,�

G�:��t,4쉎d֏рE�-P��L�/�P΀��e<q�c��I�e�\;�渔iB�����2�����%
E��}�ST2���~=���/՛.b�E2�>��h���::�.��FP
���+\�u�YP��v �]��\\3�WC�*ԥ�wHr���eq�Q�͢����'7r���/S�Ӫ�1j�ۘd���pyV�z�鐄�=c���٧Wi��D�ɍ�O�Z��#�G�����.��@,]�zY�=/��G	�6 >_d����Rs+.IiR�A0��e�ߠ�,W�������z����y�ga:Q��[���;
�S�?��8C��e��B����E�$5� ����p�X����ƿ����9(�x�;!�f���D�v�%P^9��#i�(Sa����W��'�;��=3c�kk��s��P������30rk4(���4��גF�ť�Y��uN+���L�<3Μ�l�S@%{x��P{����]4"��('�=�$d�4�烙���W�*�}�����<���{
r���{i�$�H��C��h�E����� .�
�UNSuf$_��W�)tf2q�W]f���$q]�A��2\<�n���&���V���
��W��SYO�1KC�)i�������I���.hb���d��z��<E�KՉ��n���M�%w(?�{�x��%�t(
1�� a���X��f���k�a�(Z=sv�ߊ�/�S�H�o�g!�a��o@ 6�� �;�5��~���d� J�M��֬� �ěʲesJj�B��/��/�㉱�����~.�^Br�F���﬉ �?��pM5��!g�:�vɚ����=�^;z�^[YqIw�O��u�A�Q�B~�l�@���(�Sm�#�j?w8H1y��@t��^QW\��x�IK
���������һ��]�:��;��&,�{���]���=m��(���
ýO���bU�=<�~�3$e,�T8��R��.���K:�uI򃄅D܃����<���Ɠ�'�-��(��aTQ:�_�7��U������F`31D�L���K�	l�oF'@��UkR�io-�����;�� lV��-	TS���,ph�<�1%�_@x.�iъa5h�eГ4;w�&�SF��U�9�kr�������������݈�z��Cz�A��2��p�鲄pe�e�i;�c{m�v�'�y[��pv"� ��F-'�e�s�d�=f�S4�7D�����*�{��E�����<���8�5$%r�7T���!Tm�1a£�j��n08ǵ�\榟<1%�~u����G�+}FߪBݻ��fԂ�� 8��HF��Kw�����������?��@�],�α9R})������2~i8@@=�a���Lawc��^+w�O�q��f�CN�lA RJn0;�9R㧷��k�kC������Z�P�2=��8�#��ϲ��12VP���\J�V\b9C�i¦�P4#�A�=��[3��0/*FAP7ޖ�?���P�\�.0�,O5B��F��h6���:C0w�@�n�])��z�iR���]���T'=������6Y¾_͇�{f��A���b�Tl���QC�4��?���@��ti�z�x�_�e�*����%m-t�������Ǯ�ϠźY#Iƪ4�`����;W�;��v�E��Zv��*u���0$i�!�<|Q{ ,0����Qܷ{z D7|�=O�����E{J�_��`�}���)���jH����1���SL~�A�@����mB���m�8����yIf(b^��XH���0-��BuC�Q�����u6SA��2�[�P�Ȫ~�^rI�Ԓ�v���o�u %mt}�����e��jL �u��������ˏ�8�+@�{H]�-#4�� ����J�j7T�v��Z�x�8�|:��u=}X���ަ�H6~�̗��1>C�V�r�4���;��f�V�rF������ {MRN�:��j��(�<.�c3	�|��I���F�������U?vU��$�!d��a%K�F�M����]p���+��!��.�g�Qa*���VT��嫨�A}FW�ԭ��T9���B�Yw�*j�݋*���لo��a�EXm�`�l���i��9�wB�X���M}q�[�3ͪ�֕n9`��?F.y�h���7��l���/��^OB� P���qM�2�5$'��'3��c��w��u���;L�?��aʓ��4� �&�i�J���>�r�?9��U�\`���vL�]83p�F����M��r�e���r�������5� ���ms=@m��,��e�a3.�e:�����(4�P��#�n�� �q��('�;��~@f@"A�ar����p�)�OBhS.�$�[M���W�4���1LD��$:����7���<L�+���;��촌���kF4i��]/���/�q�TL���|&,V��6�O���bO�k�Kۜ���E�7A�����A�3]Fj{��6W���LP�i���ؾF3uD�p���Wna����C��~Z���=�Ʊ�U\���6W�J�`DN�Dmġb���M���d�YQzp�9F�Nn�A�i8����Q�<ӅÍ�|l!_��J4�"{�~z+S~��a�7B�B���u2�?CG�-��v�8k��s:��^���7���zV�s�G�;d�Hr7N����Y�DM�`2Q�����~Y]w g �\_�f�ΰ���Y�o����YVN�:�~�<��L�6z7�gS�����S9�#��c�-r��9��K-�*xH�c��#~�%O~]A�Hi��į����n�Su��/��C�G�xo,<�'k�WO�1�%w[~Q'&m7�-���c�b�r��״�BU׆�v�5�������c [qX�x���^M�Ժ�t�G���؟��DΩ����"x�3���.����תы<,�JM�� U�OW�-�$};nH�7���!�+�Ui5����t��h���0�+��WþqN��@���E��#3�V�M�R�s)�,2U�^���ȼ�Q���݌��=~R�� �	*"\
��7���	kwTuz��5����\l��5�:,�#\&΍0�<���x��A���� sr�X|P'�@bk7u��:�����p����	iɲR���[~�B�E�f�0y�*A�HJ��i��eTw��^]
e�Pb�SȞ2�0~:y ��C�`��f��q�2��Y�~@�3�	[��������gЉ�X?j��\+�M��+���!A��rH~��8f�'B9�q1|����|��~LuAl.�>�:�y���2~D�sF�8�E.�]�4�P��`���#!K���Dx����7��_%�bJ�.T�'����D퍼����;st��.l�������i��k'����!�����VF5�}�N�U!VV�]��>�l���\��g��E��wil�'��ȥ��/���sb�Ҝ2$�_��#=&��[�SH�84R-Q���ܔG@�ȱF\� Sz��.\Ʌ
�@�掴hk�z1��8�>工4_�\{}[shCF��905S�&=���G���d��	
t\��wX�#<�pmm�kz"l�r>Y�����ӊAh��e�ge8B�+�(pkO�j�CѲ��e
���_���ϗ������1��(�()"Ը���ߡ�L(̹"7\_j���֗+E _�^؁A"{�4;:���rW`���D'�0L��O�?�H�1T��[�(�mP��}BjѠ�P���4����O�*����l����Ö��]q,?��h6,���ߢ�Q�m�5m�����&��5�7�"�B��4s$�vj�ꠄE� >���������%f�5!�va�0$jڸ���Ԉc�����Wʑ�B��5'�[R�+u����R���~� �Tm88=+�n����/w߼��|�H�d��]��r�"{�)��)����q&��&x���`=E�=��Cg�fx�� }���L�6��$绱�f4d'2xտM6��yZ�kV!�mN�ḒUˮ=̦i=��F_�r�kr������K��z�Q�R�=7�oSk��ѩV��v��C�h��J
M���ӄTd�TD�l&8m�%}���,�a 6�s&�$s�F�rR;� Q�'��j��Ym������gseq&ϙ�ףI�Ir_g��vŉ]�̨��-�������J�D���L���y��q�e�dꠏ$p�?l2@U�x�����]hlbn��u���LA��LEw΄>�S�ي�Y$N֍J����'��}���b�r螛����v�D�C�m�7����#���ZFb8	C�H�}_+!�Б����E�+�S@�ߡ~�IVW�jHi�ъ7��#@t1��ڒ�[�VO���	�ϚQh*�� И{:@��YF�����P�B�.+o�E\�:s��qS&���e�O7���k#w?�K�(*��Q����{���8�My��������?��X��0~�+̌�so��$:%��N�숢�S���4ڃ~/Wы�d̓�*S���s5��v�d��i���G�/$�1b2�A��4C8�fIFR��W)ߧ?3��Ys��C>Ks���t�*��]�`ӨF�m����Yy�c�&�6���@t�ݪI=�p}}7nf7�\����Z>��9ha�|��?�K�B
Ł�L�x�O�C�_[����t:3�n���P/r������N'�yxO;��v�-TG4�z%Vv���;�,���^7A%�r���v,}�/�3����z��ZȪ��x���cr~�Y-c�Hgx�!+_��;d-i�&�1�M@Z�5if������`���iG�J�I.��SF���(ՠ�2��%���Nߎ����M�'���Z_�V���1Fhs�;r� s��`?إ�M+��`���F+��]�����2<�q��n�o�^�ݧK�� ~���e�3�������U���К|��"_O=���GȮ���0�_��d��L|����e�|�NX� U���-�c+�����L�ĕ��yR�J�sԟ�� ʺ����x�!~�Dg�\1f���;Jl��٨��%�wCz�^"�}/)�m. �d�/1P��A���b�U�Sdᮿc�-�֋��9pAH�ã�d[�p�{0����q��<�j�_�)S�:s)��s/�yO�J,v�q�:��F�L�5�͢gs��'�N�L�|X����*��qaY�̊��
_$@��?�(� ��5s�6������B�5-�[tmF�����t����&���f�$�/	����%J2��&#�f�c��w_j����?���I]x�)�����f�U�h2��`���h��\ LP���I�s��a\��E�����^�b AR��o��a���Be���Ol7������"<��\Q�Qg�܍�Hb:���/��Z��`���'#U�xj`�MkS�H������-�/W�߮u�j���Eh=X�Q�d�	�h�w]��C�bD�qm����FL��q54S��'�'T�^�OK��9r�"&><���b��D}�w,�_-�P�4�(��
�{�$w?)f�i�[A��D��>(�£c�'����c���>��܇��٫�g%�9L=
�?\�)	�ȗ8�Kf�@Шh1�G��]�A�I��ǒ�|fU@��O��l�i쓌�Z)܀�z-����k�ee��5�S��nIʑHfSJ����u��!�-���}/��vo<T7M{��ŧF�U��H��Z���}��!����ݦb��%ѫp	���k��)��Ӂx`�Hև��T���c���^��xa���'_6G�h�f���h�؊;y��V
�Q�Cۜ�a�6��;�@V�!���bD�32�(�IwB��D��!ġ��]�E��moY�G�;aݟHP] ���@�Ӫ�����h���}�|��Nab4�dT<	��j�~�pWGj:�/��ks�F"�g���$�MM7M�j�M����:Y�R�rU�p�Fr+=�p�~0�\C��{�z��!��t�%�-�����(?2�ͣk�ٱ���l�ג���Nk�P h1J�l���7�u��h2�"��=��Y�uPl�U�XlxVHYEB    fa00    6ea0gsy}TH6���}���<}t�#���)2���g����M
�/W�lipĜUX_��)�	��%��8C��X.w;U��&�C�x��R���ϽC�B6d�yV;�J���x��~�ܹ��W|�n}Ⱦhɴ����X���M����]mm0V"����i �X�\6��k2��t��C_a��;8�y*����%�F��V�q���k����-r}yP�U%8*״����*׾!��_^'��#��Х#�Z��� uI'�a�U_r�9M\Ңo�NI�/�tO3LG|y���i6HA�yf�BY{�и#+���0�b4���nP��-i�� �&]c5ސ�	���*_\<Ҏ��EZ�P�Ȋ�.bE�9x����+��R�����6�F���\m�_����Kα��Mv�J�� �w��#��sH��<��f�����������3)t���\;*��uJ5N�$y���錇�_����V3B7E�Ը�t��z�F���`h���N��f�5@x��:�Hˏ�щS=j�_��v|^PgB�l�͙:��g`�%����ǥ��GL��C(-����9���@��Y8�3��9���r1
��=��f	�H|����'�ꪔ���k`ۉ�͏��Y����Y����r���@����r�ٵP�������f�<:_̭5������k���Y�pc�
�@�Ӡx&I�*<�lbu��:�����S@�b����`�*��X�ᯃ�t�4��r'2
���<oAo^�� ���P.�]�s���~4�����b�ܹ�~�2`�(3/fn����V9�K���0	K��9���6��ع�9�%Ҿ��v��,B��.%��u�cx�TZ���Ɉ�K�.@�L�y��0� i�TS��bZ�Є_��4u�Z�+Z&fw\�F�mf2 ��C~���	�-�1�#�:����L��2s�BG�p�@�2�6�A�76K{e�v#�B�Z]��T��'V���m�e9�۫��S��z��gq�(�8HU*��{��)����Ja&�~ǜ-O�C6�R�xr�����?HJT(_ý�ER��֝�v��z5/���`�ۓ[kaB9�����uG�Q.���Yc���^gG�j�&)  8t��YLM��\[�}��=T���rD�^���6�y��1�X�{⃈�l���vdD?n*��m���xٶ:ò4\���	�˕HZ���3~+A�A@��ʳY�[����/����e��B�xw!�t��h��A�YMfmd�e
z�v$0ɩ��-�$�Tr` �V\� T�%Jr�"��u��������f��l*����۷�=��2��b�Qt4� ��}_3���v�ä�#������9�:���,d殽 |�m�,�?���U��M��
��N�~�
4�%��/\��s�nKͺ�t�h4�uQ��n�1�å�l���L��z4��f�4�F�M�7+KY�u"�>��%��A��6F� �B�1�^��1�dK`�T����=���k�ԍ�m���9W��f8aަ�� ����SUV*c*W�R6�1-�l���B��E���t,?�.��e��o�"�q0����_��Ή�T����s�ը ��������~+����J��WY�ddw���w]^����.��sC��ؠ&t��]q숰X���eB�� w('��t�?��Hg$%�P,B�H.p�#$*7����N�J+fɨ��M璞}9�k�9'�X��]��
��e��.oE��apM%�BOP��o����"��PV{�7��!P����;���i~���� ��P#S�2��kiU �޹.��˰%�KS�Cc�w�͎���4�������br��Z���#��l�x_T��B��(��۞x�cP42u$���K������T�o(� �Y�p��7N�V����I�C(X�=x�����+��麕ԃPKt���DW��z1�R9�V�<��A`FïG_6S\_�;�\�|�S|�:�-���Y�Xȋ2��~��őr��i=�i(�~B�a���P'��	�W-���#�8����7����ED�+$�΢3�M����&�Z�ŗ���n��}�F�=-�T���� .�瞊�̈6��F6T_�@�y�����"T �k��9SN�NfRP���D ����+�3'쒓=��f��������%u�([=�}��y'1������/�o�^H�һL�U�I=���pHohwM���䀣��.�ƾ�Ą�Y�JHU���-_5%?讒�c���7+j#�rN��K���*Ja��������F?,�+�$�%�t�)�ng&�+7.߂�E[RI��/�4�;�I���[6��i����i���aC�����Ҫ�����1NI��姺���\o��t;�]�� �x�k}[����B��|.��møH�!=J�ț�q��G�v�nP�~����������>�!�bq1V2 )����C��z�x�$$L��;��硾Ce���C�C:���R��W�S'����I���1ߖ�>�����{���ǎ�!r����m� ��kxv-A��]��J�q�.��FG���IIֲ�*��b@��cg�ڝ�(v�J¦��DK��q�c%cf9���?���@Q��_�rq駰T_�%�^���,)E1�۠�!��v}�O�s�ٰW�=O����!�/����,F=l��U ^�e�h^� �E��ꖜO)�$D����l���V�H�c�9A\���l�=��b�\Q�FF�~�);7�+UF����^P�)J��Yg���>T���qZ�=P����{j*�L�H��8W�����7gU��	���d�'����>�:��;��JyB��2P(ݔal���%C��"aӺ�fAL�����+u42��c��_��u"�a��/o��A�.o0�&��nߦ(��VciQ��R�o:�g�#���G� �9��*��U�h �e �IIF�-�BD~��)�֡G/@�-I�V�%��B�QX�^��n�OT�����q��p���S����M�L�� �U�m&���ݦ�AZZ�v
���u�Yl�-g�h�_�xZ#�&v[:�c4G� �j}rIG��y���?�U�X�\kƣ����A�V^�!T���>够 ���L`� l5Q�.+��Dx�5���L �S���ģ����JN��I_�g������yW�ヵ3T��q��v�~N�wZ�`\�X����f�r��=��f5���l�[�&e���E ��f]Y4;�ڠ���+9����s� wl�\��l(�mB���"P��6���ɝu;m+�-I������Ĵ�?r����TzX��S��c"�;_�������o��Ȏ�n`$�q���D����$?��"�۰L�8�]z>�r���,,α�]����d��HXG��ǐ;��-
H:c��2��u�}bp�ȝ}wI�˰��ym6',G	@�<񘏄Ӟ����J��I���B%���K",��d�?`�>���i4K0�,����B��ݽs��N����������U`(�Q�e�������>N�.�0���7�7����O���R���s]�OH%2�|5ߨ%(���l?N���yVK`�2Ƿ�K��������qbJL!q�BYx��M���5�7Áeh����T5�(h/\���3��B�1��ߡ��~3�G��V	bf5/�~+>y��x��/�����C������<�q,(B�ƒ���e���eh�5Y���b���b[p�.zԕ��ދ��|�F��XH�d�i�Ϟ�o��_�V>�8n�6����+�n)
��o��;�Qe��f��ږ�k�&������(�ث+^?��S���|��2�	�W�S�Jf���y����Z>�����S�pSt�$���G#F�z���6F��f����?B�I��&��f�����P�'_����;�U����S����X<�[�m�7�����O�륺 ��1��w��7$�U��!�x���1?�.��c T���ߝl/2��L ��n��?���Wg�ţ꧊�N4(����1�I��QRS��=]5������9��$̣�ͩ���|��τf`��O���q@ň�����d3��Hl6����2�?}���_∱FHf�f�����9]��񢉿?U*6�Nk]ӛ�dY������r���M|��%�=��s��l�į+z�'Ւ�)�������U��Uo�ŉ5���yV���/�j9�[�M����^>ST^�	��'k`Fϐ���t͘��Z�ډ��3+�3{��}���ك������D[�'���r{%�2`�ݐ�� �Qh�aW	���ˇ���nĪ�;:s�ݟe`t��
?�C�#�Puu�����20��hk	6w!�,�$^�L,�K�.l��#-a��^,��~[�)�f1v+T�!^��қ(���lv�:dtSv�69]�o�L��bAj�hO��"�d�n�B���kg���N���-�O	>��	��������@������&� ��0�Z�ڵ �\���{`�EyBU��]��@>%�ǂ�����=D��o֍-o��6�3��"�N�F�Ly����?l�l!���.���`+�̇��=�`�;��W��M�_�K� h8H�������*\O�~�H���Cб�f0<��_�(	�V�Ǯ���a�07���(��ݍ��#rz���l"��$�M��(Yy� f���4%֣}L�ɹH����o?�1iě9!��"�7�I:�L����Ɔ��=ft5�̄���,_P�Iǹ��&��87n\u�?��#e��=B�2��.�H���/j{J��A��f��P0A�?��7�.�F��q�%�v��v8b�"�!�/!�\�ֆ�̅�Jk��:/����Ee����>�'F@/lv8��5�組�����G �fjd��}�>54n�O�8�6C�G}V���e���h�'��uP
�F.B�bTS���z�O�0�K6�(���7�z5ҩ��NwxRBj&���G^�%	oxx���PEv�g������с	l����u��Ef�q�:�琳CKv����q�MH�◞�߫6:Y����vr�3�棭��f_�V9��	�1��N�Vi�ݳ��-�|��������L��x�Z(�B���_���JS��6�(���K��\}6ƙ��?���:�" �Z��O�7��?�B�Q�������,��S�5C��YWy%D'�z Lo�-;��2���R�I�ei�	�9������6X���g����r%r:�G=������*	����*}����f��ix���x��gOf> Mڴ^zĩm��������T��>��h��_]���,I��O2�hB[��.n:��M�e?��]x?�������o�=�c����!�<ut����=��?��{k��@�豂3�����zד��c��ԅc}��ު�������.R�?���G��b��1""c��,�j��f�i�B�Q]�Z;��g�WF�? �_���:�(���#�dv�����D������:�|�L�YU�^_���Y��$�G�>~�Rw�0S��:cM�;>��!������*�]��p���-�� V��m�#봀������لZ���������͏ٟ^"
������X|��F���D��	�
�I��:��>D�p@1 ��w�DZ0&����c�?�eO/���.N����c�$���8�8���zufw��j!�{�j���̪K���,?����������c����_4��@�Ѣ��^�T��w�	�0E��=�]`��2��7]�u�E���:��A���Ӥ#������
G��<f��Z^��>��_({v{ҧ՗/Qa(���v��Ĵ<�m���t�EB�����B�8��աc��悢ʬ�O�!ųmrz� c��&��(����r'?���ĕ{��ʺ���zk�_i�Sf��,�0�TT�G�B=k�mc����K��O�3~��r����*Lf��(�`ʞ�e�EQ&.��Q1�]�L6\���k��2��/W9�}UDs��fT%q�ds&C���%#8r\�Y�*+QF�q�Ŏ�$O��X}DP�iK\*��m�Z�4� y�k ���%��-)[]D-���Y��̀w�l�Gf����#+��w�m�>Kl�]�?ݞ|Y|�����s�Vӣ�V��^�ɡ�g����6;�"YFl��IM�7��~2�P����� A�6�9���f^#lg��[w���|�dM�n1��~Sn$�D�1fh7 [C��b��y͇��u��v�{T�R {�Wb@��o�j�U �R�@q̷�lW���SP���͂�N�!�;"Cw;Qp�T�O�ڄ<:���D(��j�(~�^�Q�|��u#�P�AE`���V��X�`뜞&��J�	��=TT��տi���nP·�kvp�E�y/���r��j<"�����?���/�Nd-]@���� =�������t\�5Åc�0#�gaI����)����ʶ}�7�|��w�#|�A���>J���V��j"��qa}x(B��y��-�~����o��n���H7�0Vp�/��C��e��-Z�(	9�291��^�����Fn|�������D����v�B����,S�g������������t�\�L(��Vx0O�`���[��#�F�r�.E�F��$<�uh>��U`�yB���/��T��"��'��Ώ�������B?�f���bn�M�Q�M�kYu�+lD�P��M(���M��` �4�C�_�� ������	rF�CN�0-�\C��7��.��T&��vua� yt��:�FJ6(k��[��a[�?���-� *
��R���
�_L�uB|�s�����ˎ=J�5�̳�����ԙX6-�N0�"7�^\�������X�ӊ?��^ڞ���&��M�")Z�.�С�c	�U�!�"y�+�,j!1h��� ��L��,�a6�|�[�C;��x.��m�)�vw.c嗄Zp�Nr�T3��m 3�@�%��?k\l�"���%A�����n{D��"pKV�D��	�����,e�z�*�ACS�&��!����{���%�M�Aje���Ԛ�gp���}[�y~��b�k���r�J�hV=��p����` XZȯ���|�/۽P<i�b=��v�1��a��S�I!���:��j�B��xֱu�L���X�.C���':]f��N�[M���_Ɲ�#܇Z�m6��_�{����j�L�rBXOa���{��}9��\.r�]��_�9]���e�l���'u~��j҇lw�f��"ޗV�e����@mL�Llj�ck*�)�,ьo�0v?+����<��9�5)i�W��C��N�xc� ќ�cj�@P/���݌e�]��2.��Yd�'�U�B�	�k����N��I�3^�+�2�C\�^�����_����(�g�@��]]nxJ�8��p�	�
�ή��m��z��;q�g�Pd��z��i9Z0�l�>O�]�K'��Mآm� t9�n}k��C�=Yu3�E���*S�=�E�%�\��`�O��]:剩�z��$�X���3Zq�����0�_򏂭��{�v��=ң_牖�2����ݹ:8�(j��1Y��l�κ�����> �I��l1<[=�%�.DAf<b�~��'�h
��5*d�}
aC(�\����8�7b�r8=��&����q4yC������-�:(Bn��<qG7ԇ�Y*�Nׄ~�Fz�T�ae�e���r�x�m����ۓ2��Њ��p.kݫ���Kc���S�o��S��
q֦���I����Vc��ЛS*�:�������
��p
���L���` Ƥ����B��:Z�z�`�?Xs�J�<ss��vH$B	τ[Δ��j{]��ϱ8iDf����qq���(�̈́��J�#�/� �.�u+<�z�q�KW�4f�]�i���I2�ձc�$=hW/z�:���|YK/Xpd�U��{4t=_#kvS08�+����ߥ^`�]<p7�VX/!-�%J"��i�(17���LD�$�
�:�}$.��:��_zbbY턮޵�#=-��Y�]�'�c�Ԫ�����b�pQ�T`T�|(�"b�3d�����fX8mV�񸗫�:Z(����b�"�С����J�6��{Q��5������Ɂܸ�-�7 �~Q�_{"���[rtZ�������훋�Q���V�W`�]���/�[?#p́�ObA��{�M0�/�r���/�0?����~`{�����*S
��Tb}w��Y�@F���{�`Ij�������+�g6>	��d�7���W��)*����!�!n@����김]P�����)u�U}�gR	 �B_j�'���~�_�!�L��3��*{0~�R���=y��i�[$An{$Qf�~ �ݦ��U'�'A琨�Ƨ(~z.�q�IP��~:QMX[�T�<�kZ�w�V1��ɳ����~��0�3C|���P�xRCcG
����d�:;Z�5���]5�MB���:��� VƱ��9 i.&���;��'�"�_��iA��4,���u���ћ�Hޗ ���Y�?�)�9���\��#$j�K��u4�5ا0y����knƿQ<���/ZO�#�lx*��B�������,Th!`�`��(�O����ӽ�`�����~N'��.L�	��9�b�U�`�c��*-���Z�p�L���r��n@���y�����]8���P�^R�gL��e	�)�E���j��;H����?�b� �Ӄ*0G��Ѯ�O���#�R�"�"ʣ�`0&V� �&���!SJ|j��q����DN���]��&� ޙ��v�l�1-{r�3�����5J���z1n&4��҄�7%g	��[�fT�<^��?��K�(ܥ�S����SL���Bfz�)<6�z���Q��!ї��Pq���d��Y�ǎ4$�?=�;\��o0�U΀���fbF�ˬqe�*���Iws�d��8PTM=�"*�zd7!�q���0����������4>����pw���SǐC����.O��Lm�yq[���)2��ç[z�;n·�;di`T���+{�;{;|I�*:"����)շ�?���b�o㮔V�@�cf�<������C�vpw�mwj3���p|��?�L�Sނ����1 Ss����i W�~9�hk�{�5�T'a��#�������B���y^��6�[�����N�U���Å�1�&��V���dO�G�;�Ƀf�e�y��+��A�{p:�Zg�A�oS�?v��ܷJ�v�T_pqM�Sy�%1�ʋ��a�xah
�
�)�7�\/����.+{ѽ#�~(v�!�!��E��E[��l4\4���I(Wki3Ctn��:q�22FC���,{�t���ꑐ��JVJ-�Ǐ� 19�0�.i���#���3"N5u������ax��k��d��� �N���d3Ho��m󉢞`�Ӥ�[�y��L���C�t'WU�grxez�<$�a!/1m����y�9-�ޔ���d3�_�����󳥐/Q^�9�ˡol��R�N�ɇ`�xeٺ�����:�P3��J�G◩hN�i��~�V���a��l��g����) ���-f�菽���Z��:�zȡm(L�)�K�i��!���x�k����n)rw2ߠ95EEf?$�֎���_a�ň+��Xig��ga�ѱ�ҭ�P��<�{C�v���V�v��Sk��Y�D��Q ſ��ո�Y��y.U�v�,zAS�j��Qv�|)Tx��a/7d扃����t�����A�-��l������w)�u��f���&��jֻg^��9Vgڪ|�hTd��o5�R`j�S��Bp�k�l <g�]b~�ȝOFT+����Q[F*HW_�*ָ؈��4L;��>m�!M�|3�EQ�z�w���5�D�)-n7bd�iyYk�<��b�z;0�C��|H��1Y���#�ϱ�p���^n��;Ї[�Մ_هD�[�^r��y �[����(�x>ϝh�,�T-��TֲZ����33œ�m�g�����`�n�r����tv}p����>!���Iw����q���cX"v�A�s��Q�Qo��G*YI�a	Ĥ/+�d������*P4��i�Re���ӱ����%��]��9�u�-m�VZ������븞����S�څF/k��[��P�h�@��)��pҀ���p��!�[[�J^_�Ǔ�ߦ����
cG�S���ZYǕ�V9�r����l�q��r�.8��ፄ�)�eש
�O���}�"t�Y^��	lk�Q���y�A�	㣮�k\R�0�U/�޳�W�����0������J2"����muk�p[]&֚�ծQ��7$�����Mǘ!�m��E<q��+����0M����tr%V���R��Ʌq~}�3�p	�z�~2]�C��ܬ9�y�]Nz�b��h��-9�R
��KlAm�*��'FQ�B��_�NO.�5ͽ~�jJ��2�pT�u��g��S�U���ec�S��m�O�Xpi�}��J�ͺ1}��i,��8h�-j�����ZSC�8-������Ö�&~ۍd�R����pM����j�QH	j��0�Ǒ���2)�|J�{�qNE(f;�%��$Ư����9 ~����XZ��|@���D�Ը��PgT` c�� *���J�j�����Y���-pɹߘ(�睟��G��$A*lIk�/��Вx��n/�?� ƥu���1p�q�m�e���j��oLd��p`�����P�T�F����A�]�Nr�� &p�+مO�T��O�1�iA��f'u�)�Pf�.�|���B���f�!~�?�� �hn8l3�h���zg����Bo6n{nD�pT-CL�4�;�I�1�m@��;�/�?�T�c�:�uP��=޽0�Pu�/Ԡ¢��t��r;�m�l��63��B��L�ٓ~��70noW\�v4��ąSY�ކeR>�6bV����Ԗg���Q�X�ڟr:v,��G���]!����_t�S��OȌ�����XН���G�WІ mΈar������$��H�bF'	F�������|��hi18��M��fB:�x�a��v�?�qx��I�s����a8�X��[�9��<Y��5L�Z��1I��&��x9V�%�A�J1�P�H��8{eh���ճ�Ϗ���2o���&�T#�ڤ�V}滔1��_:�u�7�Kk�V�ؑ�����q M#�6����AXT�g�	�roh&�̥ �n���L���.�S���S��I~&!hp�E�t�Kw0�]s��05""�q�w���*�^��
��r��*'�q��6����{w����#�u>����Ԃ3s*�(���;�(H�aPU8o���1��F�@d�̲���x$ap�<��K�ʱQ��n�����qA�s#q��7�#��1��A�l�c�E3�*����������ғ�S����x����ZQT�d�F��-�h:�5��(��\?O�P)5s(��m�ͼ�ibI`<��Sw ��Q�3��Ϻn��q%#I4���:=]�Ƌʸ���ħ{1�ćk\��_�Mk-B�$�Y��<R4����=n!����VŗUϚ�7gk6��H��XgE?�aA�Q	�8j��l�b�UACb5��!#��>d}�~!�ږ����K`Qs�lc�����rD�Dp�F؋9���}?��Y��EYօ�@]H���4�S������ơ' $i�>(�ſX�ǖ����7ɏ�!���v)�{�g��Ї���w�Ԗw}&��T2Ѱ.��^�\��U�
�Ԉ��~e�h�K9��4���T'x��^�V	���Ȟ�ɓ��g]��:�b9r/�%��68w�]���s-A�����$��a�b�@6ŮI���Q�S���&�:�� �8p��K��GV��T$�?n���%KHq�X�tU3�9щլ�Kd�~q0Ž�<Z�����ȑy=�ϼ�IɶS'��Z�0�vd�bCזUf�����oP̉�����ji"�C�%��Юi4 ���>�7?�0#��#ӆ�׆�ɳcq������@�S��׃���Bn8fn)�B���t��I��eQF��X?j*�Ŕ���X�-M������e�X|x�]�a��m&�žrT4����{�t�Q;��[���sz�Yck��l�]MT���h��J�N�ni�����7KM����.��ƬP����)�g㘝MkLm/��N	�*>�~�m�W�t�X�}[5����r�Ԟ[зe;�J����������{�Qs�n)D��j�>���:X�\�p��ԋ�l��
=T#R�&�w������4�ߤ�2��]������xxAlR���/dNn����AP�1q��2G�v�(��2.J�e7ם���E�Bx}��SQ�������ډ����>?9�8td#3$��hS2+���A��T���>�`qBN"�Y����$�SDyM� �S~��U��5C࢈$_2���AL�F�����#8{O���\Wm�N�o�ݎ�/I\��{�ߖ�¶^/�U�X?T6���|����`?i�ь�V�L3�	��G%>>Ї���<����V±�����z���nJV:�:�js����;̊�����AV='p��%aeˉy��+:e��|�9�x}�����?�H�=����Za��Yd��:�D��(�.�)c/IU=�(�<�L�ZہW�� ���fsO71+?�,E�䌗8��kD��W��3U:ކ�B7���g�w�O�"� T�Q�Kld>����X���p����=�Lk��ͅ��"'@�k���pPFłܹ��P2zn�cN�Ϯ��穌u-iyusx+�G�ΰ�����Nv�V�8���>VM�v��ݸÍ�-����W�������S?�2)[�77����kmVsP�l��`v�[�J��%��z��=��u���A�e#���Fu���pA �Wb���ʌ�m!d$~�����>��9���}�9|��'���7˹J��w)ka�Go�A� ��uP��4�Jŗu.|K;
������7�]j{�����k�6"-&L�P���Krt�|�+V
�^&��䷷����%Of|�>�<%�'�lE�֗�%'|�7C�H��u��.����$Mp�˄9�C$1U��#�E|�]��f?S�z�m�d!"�}�� �.]�u�5�p��R{��}|2V���r�IIT�(�P�d"la��7Y�e!J9Lٸ��7������X���e����(�|n��V8k��cY�n;s�k����zh)g����Q�.�H.��4��et����������;: X�-���:�|����$'y#V9�)��3��I����x+�v��
���GPr0�����>�_��n���+�h<�й=g�=����$��_��Ǿ�M>(�J2���d2�[���~�.Qi˹���/��j�0����4+B>�}�x̯�a��3ST�����/f�p���i� ��A�aU��fA�x�r 8s]}�VV����n�X,�#@���b�ByL���g��.��v���w$8"�y�%�\{&�u�MB�ͧ�%^��K� �I�MP6+�¯!�U�Ԫ�M�x��g�Aq0�!PF+GϤdr�L�f��9�����pՠ
'�t��Ì��x��B�I��0/��q�i���\1��,�#򙮦�Y�'b���Ys@*���u�6�q�-��\z�
(�?��Q-oTG�O]ܝ�����0�䰉�[�$"���ʞc_�
]����j���R�w&�WY&Ŷ��%���4�'�Jb����Z����]&k�#�IH2� !I�{����~h���q&�D�?0�����=��q'�4bM=B�T�̶c��]B�~�řP��}�/{a�dѠ�E��j��1)?)�|�_��6�WI����ޒ3��1N<x���
�����=P��
Ί�sbٳ2��m��"k;�7�j��c���^�y)T��W��C1�/����� >#3%�����Έ��,ֽD���c��*B�0q^�Z��q.������,�F7u�=�β�ڭ�0�fɘ(������Y[���!7��\����
`�$�a\�����u)6�M��3�Ė,0;�cɀy�ژ"�>S� l�܄Jh���
��شS��g%~�v+V�����W�d`%"� ލ[[*	v��>�������-��LvTW�*-?9�@{y������&�H�����V�i&=�����1�9
�F�@B\Ϻ�8J��=�$�\&����t��@S��B��I���~��n�^�r`�G�R�.�&F���*���+�dK+{�O�ouۋ$��,�����w���Ϧ���b�b��v5��X^-���Yo�+�����U�㶁�#���ݘͅyъZ!� �#Ff�V��]��]���$R>/�m�'�$I<#m��.u�fj�ޑ*����vk��N���O��M��R��!���,��ߛ�C�@k���HT�q|[���_�y�%ѵa~���݃�?���4�����cC���q���̏�O���[�i
0,N&5�]$M��"��W/��^	��)q`��tA��/� 	�e�Zݘ�����5H*zT���Y��O�YI���۱��N���B����^,6��d? B6�����MH���tp(+�OpWTr�_֤��pH�d���4*Y�0��x��}�	'�j�WL�|j�KXd��I4�KLb��H��s�X�$�y�	�G��Y����:��������B$�z&�ʟ�r�����X�g� ����� 5�cA��]����^>f�P�s'Qܤ~�=KE\w����R�������N�����|[��f�����e�,BrU�=����v7������g���W�ѭ�T h�&j�/��󍶻4L��釬�8'���Ѝ�Q�]�A���olC�Ȓ��N���xr��p|��>���H��E*!�v�n�)@ql$x>��{�KN��_��y�^`�A��X��)j<���aU[�Z��)A�����T��4�{1��m��t�n���r��/0�@�懰s���8��%�5�0�ĸL*U��HU�Მ-|q������5�Ey� � ���Q��7�p5��+9ޑG�3�>��5�bp1�B^*�,�" /�� ��|��X��I�����T����v��8ʋ]k�%��s�����e��R��FU+�LV����<���#�(��-h �%EX�i ��y����)�5g)\�PG|���>�N�ժ	���e��7�2O�$�0��M�Kh?�I?�vn*�}��-���XI:j��ç��g20ҏ7?իڥ�t	S�Cáh�oۍ�3��1)x����Ql��;]mXW�)�Y�}t��U��w���tD���qD�u���`7YKy�fA�4�*�1��s��In���^�ߑ�@խ8�{ޤ��z�� C�,_6�Z1v�EĲ"
�Y�|w%�� -d9>+U:y6�tu���5QN'ѲXɩ�a�ٺZ߻��l�?Y�N,V<_ľ;���8�x���:X6b��^�������g�T\qX�e�5�>�"���� \�)3ʦZ�Y���1�r��"�&b�syBD��<�Y4u=QG�X'�0d�Zio.7���iry��o�1��T<T��}P�Y�b2�����_�=���)�Rn��*�������,�[��"%:r�|�E=s���]�C�/����gd��e�r~6�)��^O�[7��@��C5�iӳ �/ ��A!��!<	�����M-�a���=4(\��57��m�@��!,�řE ��Ȁ�u�>,Y-캀�b����_���6ߖrC�R��Xj��n&k�L"���;+J�C4\�c�Q��1~?(A�Xǩ��|��U�4��B��C/$�ɧ_�O����"���ŲC�X�v�`m��MW0yr��yՖ���\U D@��AE�3G������7�J&g�O�;BA0����OݵN��뱏�bpJ�� �Py!�b��z7�	���eG��@9M8��R����?�+�E+�秉�p
*G��]�{LCG�-�M�"O�YY���B0wP�!N���������d��P	��TJ`�g6�/��0���J����mB��&�oSw�wf#a�b�/���>�,� ���W����i�#H~z��r�RJ���b?��n��]vdۗ,��x�ɖu�Ǯ��QZe��e�Ze��[��O�r��X2�����*��n��oF���2?nJ�l����W8�V�h�Q������������-4��+�|�B�o9��N��<�9�X���!
��0��th{���� �x���[@H���%��~�Ajx�.��'�ء�4ﬨ3�4���T��l�5��p����o"��J]H�����ٿQ1x�!����zsn�s�vp��D�����#p4�%�� n�Ǳ��1��(F1s(��� �g�*,)HE�n�(��Fض�U �S-����q[�Y�*����ݵ�v�|�~�^����s]��L!ctO7�?e$@>$bѧ���k�s�|�M�o�J�EK�}�K9&��5B�T1:\�Oօ���_�;�[N�x0����K���o��xb��  E;K���΂	[2�0݉(c���N��/��lZD ?���������\!a-/��|	����^��6�xY��$ų���N'<XJF�R�B � .2ѷ�0����Q�=|H�N�.�_s6k<�����o+W�!uEy�6ޘG�o�#��H�k]r���K���I�C���m���EL��6�eo������%x�fc��!m$�1���}��[sf�a���G��a���~L@C�D��Z_��P;+@�ZF*�4U��D�\p�Iu)ڼ�U+˩ዑ��?�E*���B�n��qN�3?:ǣ3#�PZPJ(��u�n��nz�^l{�T5:O僘Lsl��a�=B�"�3�$9U����㤑E`j��jfP�Ľv��BN�/����I�P8�&�!8�BG.�_��F;���D�רU<ű­�pMF/�
4x�A|=����O���A����hN<@Y �7p���	oS��`��_�#S�i�wQ���Y����T���_�E4K�F-�?RmZ��u�H�]�#o�7���8I��eZ%lV
`*��#o���zM�ڤu]��"-�m1C�pL=/�r���]���x� �U�l�vD
��rl@�����	�jh�l����N`���WqZy1��,���%̤ҳmF�ܺF'i���HEjk�T�}R�=E��7Q �a�_�3=4h�T�NV�3���O�$
eȸ�J4�^y�!"�3����n�C�s(
	�qv�w$>Rq6�9�����X `�O����I&a����nt��Q]E��ط�`$��,#)���C�k�#"p�iը"�=��W���d�i��+U��D��(�_�r��Ck4q,�eA=����\h���0��A�یw��	�!*�[!��L:,�l(R/�#oydH]/��B.�������2s��������5�=�9����kX�or=��MUX��.���@�e���I�?�Sl�°��"	Z�g ��'�c�|��yHlS��t�v_�!�������l�um\�^y[����X�Ngx0�l!G���iuJ�!�	��_��\���l����<;+n���ƾ-��1�+	�9�.�zF�|�u~+�v!�� �����>��E����+˳o6�d���կ�t�)�EsWmި/����+)��9Q���j���S�3����Yf�;`*1N!ʪ|׫�g�{r��u�㶒��g��G�J��F�\��a����@z{����U��0O=���Q�vh��	�p�2@��1�no&N��?.�5V�L�`h�����G����
�.�s�۞ٴ�%N�ϹDb8]WzB~l��=����6c�j���#��:{�;TZ�\b�_��b7��;�G�!�7e��r�".��̦�T��28�D?y���&��h��� �)�|�ܾ�$K���HcLlo(�����.�l#:�̏a�y�|����)��K�K;�\����1~js!�+�/@>@�9��\渵d�����r� лUNo��Ҷ�ۯ����ܜ.yM9ˀ��3����~�
LΫ�ǂ��/��.�9H��ۧb��ՏlΈ����n�φ�u��9�T��2���h��bϯ����!@7��*��<r)=	�cTt�Ă'KbH��*�����*�{Q���>ȩD�G}(�d�j	D��dqY�v���d����΁_���m��A����L��%zeJ��Y���${�c<����Y	 ��~�w�؃#6�5#�@<*�}8���5bY��u�P�RE*�����4iuh,��-�(���;�������d���mK�T>�z���G�vBZ��/C��6F�-7oPfu��c��洜���3�մ�.�ɯ��1|����+�,q����i�×�RZ� �>I�;g��t�²{xj��ulo�1B���N=fW�mA�n���>��r\8��M���c=	J8-���RA�Q�����^���e�@�Ā�c�W �n�%k
>F�g/�_��T��i�fe6���g�*�+wF$~PaN�l�%P���({7�j:B�:#1�r�6�~=���>%�ƸO:𢠛s&֋D�Z����-��=���K�S�(�*NV�m�3I{��SQ��{A��Xt��7��rl%���<�3��������9��F�۲���P:��#.��*��I|���ޘ�T$q��(e�{Be��|�j?4��dИ݄�"�55�+ly�\��c��9���`/�	����r/�X����/&���)�4țsLZ͘�Np�9[*�G�{$]�^xx�KRs�ۂ���(ٷ��T�M�FiC��<�0��6���@��J���Rs޸��6����C��ux'+���e��D��7�ΆC(�Cb�L`�����ph�����v	3 `S������Y������ۜދUl�2��X'�\��~��^�֭ny��Xi���4�ڬ�Ndj� �h5}��o�4pT�\C@oe��+pe����iΙI{��?}���qµ�p��&xӥ�/��-�N L�#�WQLO|�Μ	9��SO��(Um;��U�u((�X���q�P̟0�,+L�\�.���~`�Z����M�D�[嬉�S!	W��O��(��88BG6�����h,����F7;Oϓ�������]�TZ�إ]�h\�7���ޯ���	;b��0x�4	�y�E7K�K��3��u�iy��u 5�o��DW!ہ��S��#6��zO�v4D�����Zڌq����A�U�9e�+n��,o�wh�k�;E��M�����/��(�P��Mx�(�x�i�1OW���!��f�r��Y�h�u�]�Yn�;;���(#\�$ ���BOE��T2�)-�sn_��LRV{JP8$�B���5g�Hr7�e_G{Ȯ(�)qfe����-H�m�"5��D�,O__�~]��H�zyɦ)"�PpH�� .��t#��qG��h��<���U�0ܡ�mUD��pp3�᷁l	 �[��|9��%;�Ÿ�]�Hg$�G��\��Fk<��2��Ϸf��o�AzF�	�V�U$��#.��l�#�n��S����	Tf�n� =��*��d���,�M��!�%�UJ'>cE��%��� k�&o���'Z�8��E��^��9�ť4���)�M5
�.��hTe��MU�8k�O`Y���#��:"< �ߏ��5��QB�0}|G�����^�2	N�G>P��D^��lDrKq>���y~��)�v��WcePY-2H��WIxX���D|' ��6�NPؽhȿ�/}�ס������ʒ�f�܏����!/��5���T�#@�j��@3�r�BRnM@�Q�3=�Q��;�D�(�GT�Cݏ�@���0�d��76����eH�cY9ƼT��rmA�{�GW�e��c�'9���3v@G�����F�y��Li�B}L��v�x��W�W�����z}j.j�vEiI|�,q�*�>�9������*�s4ʔ.]p5�4�H7�:�y��lZ�${<�t���O�j�{�-�cy�uK{L� ����q�ï�s2�%��J2���~�Q�9��Lk9Ia�3�⇓��R�M���,��8uD�:k�-l��o�5�D��҂����A�Y�9������8�߮[hG�
3�*"���D[��R�����Q&��X2m�r�� E@�U��'�'P��]2��f6#���	�\�፲�\��[�m��I��2h���CG�/��m��(�^���[�D ��qh�X��Ҭ�\��'\�l>�e��Ē+K��,��.6 ��L�ZQAD�TȔN������[:6ӡ��<�Gu">� �� }�ߥ�L�������D��H`h�5)��Ƌs���z�����|)�T��jW�ş��O�����q�.���w�5֓�iX�\�_�LV6��j�L����iVm2�(�H@;�m�!t{L��:��1�A7���{�Q�����-D�w���@k�Q�f�!���JY������?l��*��$=wT�:���/�8$���р�C`&*�5���u�1��0aՓwlh�`�C�����
q��6�:��E8cD��)�h����a�Δ`gq��\����+db.��$�J��mgMpd��P#0�	E]�p\(����]�ZL2��b֮��Sz���b��]��Uj���e��({1m��Q��kH�@�����J%������G"-N.7�*��uD [S�����y�f!�
.��a�:�G)�2)�`q̵���z���J�\t,S�Vy}��o��Jh��JmQĿ?1	����i$�$W��>��"���O*K'��&��W�M�G�����I��;&������ú0q�FDݑ���SFg�N
X��	�s�Y׍%��~�b�lК���u�x��i�z��(V+�J8��bwiI��VN�6܀HV� ��u���9m��y.�~����SI.г�F\�����o\�mF,m��.@Z{�������=��ax\��M��$����|��k�e��OZ�]�"e���ٛץ�P��;�o�w�/��Șo��\6T�Zl�O-�4�_zblԤ9�:�kt��(	ĜvƘ3�T�����h_,@�ut�I#`{� z����'RL��*�=����C�I�H3���_���Ͱ�v�k�<<����.)��Ͷ}�N�)��j�PX�ٳ��y(��/EA�vH8�3S���Xq�Q;\�4~ ia��MC�+�)-1�dA�Xlg]��Y�1�o睉�I��D�"���!�j��Y(�� D������_���}k>��|w �B�"����0��"vP���5Z�����H�*�A^8��?�;U�
Ό���M������2��ÅT�
�<��()�f����&�X����Ub?��f{.8p�'x��dC���x:�����9��f�U%ג�W�k\����9&���P���5�(z\� �B�k��d8#�n���~}�1���A�w���Y�i��>)��*(�:L#����1^� vTu^���1l�e���ٻ���fb-7R�?#�C�����v���_��{�Ƣ�h���¤�+Z2�.&<ьA@W �<�_!ڽs]�k#!2���JrL���m�7C
]��1�s��<�'�o�͟iLL[>e����\���0��W���"�6�^=@F�b�i�����}��fJ���T �6R��;�x`�>�z!�Z�-Y5�Ǥ���~�Nx0#Ʊ�T��s�y5�O���I�� �5�-�5�|xn~.�!$�uQ�4�����س�Z�F�p��!���󃺒鯉�@]�F�T�T4y
 �K��F&���>2\)�^op���S�H]9��W	׆⧂�q!�zч��7.����J��@;k�Q�������|�Tt�DF��J�GIs�G�p
P3�d��#�;̈���p9�	�QJ�u��k���� w��T�cz݅d�TVgz"�P.�TX��n��[���#�g�rC+C�#^;��4td���ITXi��7 ���I��<�SHj�fJ>�܉�p�m��ղ�rIXʉ�y?Ί��*��&��/G�>��[ނ�@O����JP�A��>_��[|9Gg���g�ۄ�Ī;69��A��<�{[��:/�%��]j��ch��,�)�LG[��^{��(>(p�7a8!<a ��_�U����G��k��}X�/0?A��A4��]c�4�u������I��q+��X�5&��P�@ڳq-����D7�����5�7�"Y�c:�jeV¼J��u���/����Fg�b��Ԃ	�|�W˅���Y�񱞊��Q}B�����\]H�*$�/���a�����gH�	�P��W�Z�]^�;���R�~A$a-��WNd=+�+����P�����F;U��RF5kL�^D�&�يn�C^��tӡSǚW�B`g����\>��Q����a����^��lY�NH?�CAi����J�\Lq�&/��Q�c�H���׃��DP'��k/�g�.�vW�>XLcdKu����Q���]����!(]�,u[3�֡�^^���M, ��[)@�$������c��v�����6��$rr�d�mD�o�)�^��186�t� �0��a���?rJ��Q��\���Y�,]M�\�
_�Ps�Wg�響�[jb�n�_pS�X|��r)1�C�19��`�w��mb�����q�`x���p8�ATƐm����tܙ,����O�z�
=}bt�����Y�:�}��Ѵ��ȁ��8������ ؤ,D��`m7��)�eiN��ɘ��.��������٠�����v�|ݩ�+�����x��������M `J�z�1��XPF1�ܥG%���V��τ�%��{���\E��b���_�|!@�_��<���*N|+����A���E���x��s�_�;��G��0Z��נm`�4�w��ˏ[;�o�=��V��+�E�-� ��Q( �@���\��c��o�2�����^��Ak�y�y��R��3$���� ����?18?��r�edA:�j��-��A�r�b͕[4>����h�Mɋ�O�$���.i�@+w�|>]�3��X�O0�ۼ[3Aဓ�2��R�QyC�L�q��jVw�a.F�*P�҂�	�\Xf���$%A�)��v��>�T���D��,��53��ѱ���	����Г#Ղ�^��J����g���u�F�������l{^�E絑���_��Qe�u*y�a�}P�
�+.p� ����kn�7�y/��K��ʶ�"
�[m�rlM �����j#`�/�=P�h��Jm��^�����ބ���z�Z�>ud�f�L��_I�aZ}�Z��#P����0�;�۔FĜ�����f	ې���Vv��"����#���4��������^���9��п��*�@��ԗ��J�^������y�B����c4��˰>�w��i`�ͰNJ y�P?1�H�=��¾��������\z@64oj{��ξ�ؗ��o�z��t����%�ni�jt��lx�h��40�U`�*�8j��|���>�<T�J�s	mPq��"�G2��ِv����$-9�L�7��^`&��6@�;���a�M ���d�d1�&��aV~��P[�s�{��z�c�&��ǥ/���g2�� �>���4��/)��P?Z5���`������и��>9+{�O�M����B e��W6^ ��}���h��}�y���
�{ �bYH����`�c��I����O˂���6�L�­\�%@xP�?�Yo����,(g�u!���-rNL���H9����r$�K�m��s�a�_��[��E� \�Y���hL8 �TD����ۊ-���}<��X��t���Kn󃭖��t�-Ɲ�-�O�
`�$
��� aA��ڲK86��,��I�|�����>$�+��(_��Rgu��N큗�z(��E��&���G��h�*��Ѡu��?��#��m�N��,��]��>�A�G�x_,�p���l�����#?Z�R$F�t2 6�˘�4�ؠ�I�r~���j�gR����錝~��^�Չ��e�(r�VA�ɮ<F=�#g�W�ʖf���v#[��"���^��E�5d�	�W�j���º�>�J#�&z^��C�R�Xq0'GH��:+�W�nb��VÖg��˜��z�E� �UJ����.�� Y̰�Ño|vWl�x�?^:���A�m=�f�b7����1���%�_`F�^�����C��z/�	��t����\b4'n���`��Z�&%N����7��^U�j(�%�v���AҌ�����M��k�o�����j2�E�t|�@ �$��<����Y��`+�����K�<Y�4	����О�����A J]�Q��<��Mw��¸Q�K�*���Q���vH��H��ͳ��Z��O�W�yתRވ��(�"���Ĕ���O^�m2�h���Io�0���-��le���#-��~.�9�_��d���NIU.���Y۶ s0>���Gs��B^e�~퍋ŋ\pz�t�Z�`��s�����G�<($Ò�d���2^ڨx�4�FȐ3:.Q�"�~�(h�"��<�B�����h�����G�@���׻�G��G)�g�F��)C}K��,���Ԩ@�L���LΕUFu�x$_�s�1��|.%8����sn3�`L+�#��~�+[�����x�!}��z�H�Dң����0E�,�MCx\�۞�E�t���"E�h��j$~��̪�L�$$fc=���-Ή�Fxy'ⴀ�])��$N�>���f;$��F�2�����},y=x��_)G�>4�R�_�=YY*+I���L0�.���:��o8d�j(K��0B�����zn�7Hz�v�̹��XD��F,}�6���-�H���`lи��'"m�ҏr��G)ϋ��.��I�-�s:����x+A�<�(�8pT�T![��H1S�h�R6��d�k��4ΘS��h��f6�N|=3�]��u� ����)׽_�y;�n�^
ʆSĬj^�:1��ݠ+V	�OHs��vun�����[GZ^�H�v�D«رnt+�(�l���PF���N0��R�]Y��]��*�>�}�LK|�"�� ��f��)�`p�v���7�}3��JGu�^���㹥��\7Ί�4�tU�s��Ko`��i��*uӡ�%]�?�1�->��&��4�J�>/P8����_�7q>�m4�c�P��B�pb�;&�����C1�c���YK�$�K.�$�&���Y��)�2#I�5�/	���G���(��b�JN�Y�7���QT;C�K���柹��ǽ��07�a��L�,fF���n��9x����k��J���^�	e��}�8�`Ff�$��`�h��tVDtޅ7���v��i
t�[~���u��V�h��C��B�W���"���'2�bS��A�&�mU5Γ�ɓ����K�/���\u�r�o3�Ğ�]�[�K9��p�.��!�y�����X5�6M���}p��$�9�o!�1�+.Q��py�M��6��-��b���4|.AH���n��{�_a;fyACͲ�qф(B�o��]:�9���ִL9|[(Y�k+m��nX΀�ȹ���!~u��ʣ���J��qĜB���DVʇ ��㘵�n%nS�y��7�fu�Ȯ%x�ׯ\�e]�'���M� l=�XBt*�p"���,0/�ݚEd���k{���Ux�E:���m�.;�%��f�Ç��r�lR��D��}���ʛ���H�&N���g;�H
"3�s��^�CfL��Hjh���3-_��e�
(;�c:���� �V�ҭ+3�:��M%�$w&���&����_�q���������q��w��
�5?��X"���7Q' ���Nz�kr{�I!����8)�
�Y�֎����b�`����N,�F@*�#o��Ctx�$&TF�y.�����Z�F��Z�
�[>gE�!�ǣ��,䭤�/@��^������&���������#�]��\-�Y%3�#`�8GDYb�XZ�!խ���k��(y�p&IV�X ��kY���}��r��KC0kV'|ƥ���t�NL��������	;z\h�J�ҋP�@�kJ���������YaO��F�k@ :�\:�A�?^����귘֛��ZY�@����H�T������zCO��ZKOlBe�e�T��t��V��h��K����b�'�A�K��~C҃bB>���%�;*��Y��-��	z���*�m>��" ��|V���53����Y}W�K�2�-�:���䚇)N3�������~���������!X��f]�I����@�W�p<��5&I _��/���Y��v�Q��xȪ�Ϗe���ͯ�*���L�ۄw��;���C���E���n����cw�rf�a8�]h�>i�m����V����\��'O�i0z��Qs���/6���2�;˦2��U������P�Ƽ�@�(na�5�[�ޣ����}�Z����WjU��{̃�q���6�
=iN��ٸ���۱�]��� \�s� ��8_��������_�FHTZ�=L$X�j˗�����<R�^��l�8XA�:�^��v=!§b���WE������/=Y'��?�J�Z�g�Z��5��l�x�)��b�����Ha�@�h�F�L����
��^��4�'��!��t��t��" ����:,�ߙ�Lj��U��\B_�H����r
�*��J�ӈ�,n?Oq�T��	���[���#�["(���!�a��Ĭ�P����:�
��7��u�a1_x[T����}��Ǭ�9-�m�_ҳr����:��q��|��t��FO�'q������W>�}���Yq��TA�@�Gϧe�m$���c�W����ES�d՟����2_�F)%f�"����:|�O*Osf�E
M��V���Y�iN;�=[Z��H��O��!.l���� �:h�4oF�-A@Ǌ�ʆI_[�j�?��^�i�鯌v ��:��1����]ZK�B���Hv�0*�����Z��h�#i@�����d~A���^
�����NL<u< o�DM͙�un1�_뛚�' VT�gp��QQME�TO:�K=8m���A+�4d���,Q/Ǔ����a��G:�i�$�����Ae�;�!1&I=�*��`a���쩋�=aRh��:�n�oX���J��0��&{$�-���R7s=�\����m�m�,�Z�%G��H�g��'�3�����(F�(����g-}�2������a��@Wk�5���u��]P#���q~/�^%
��5��1��)�ν��K�� �8�%/�M�|	�������I"�՚#و���GU]c�B�u��mz��­�G�z�*����Y>F}�2�^������H��A�`�%�S�)�@a�����C}�ƥ�Fjr�V}���OΪJ���(�BS�u��o���y!���oPx�k�q��f�d]��¡�y�B:
�f�dmxk@H�S��XlxVHYEB    fa00    6e30��U(���^&R���=^WE�����3H�Ѡ�W)�������W�#��Bw�\�4�d�j�bG�qf(�*^�њ���F����e�ކ�5R�6|0I�Ʉ;>��:�������c%o�Qv]�7�m�X�և���d��Z���������}��sՊU�9�ӕA?P"�l��f��etz����PΪ�|�V�, ���!m�`�����A��̈́ޫ��r��+	��ӈgD��x�1&�A�F�H�a!�3p'"�oG�T�^��~���Xt����BTE��7!��Y�kn���6|��p�/������)�m�3M/�?٘�Qz��;�-� �Dh�ȁC|�|���>��ސ��x�VM�Y@�fӏ�X{�(�c(����iP3Y���3`�f�:k#�"[)�����s�,t�����ф�ٶ/�v�Ԟj�Z���
���<�_�l�Y��{{��l�i��������&����W��R]\�R�(�!To�4*ah�H��O\$E�>2��GG����#��,�*b�JS�9�k��QA��k���
)Y{��W�s�eK��S4C]N��+�ٕ̬� ���1�*.��;:og���g� �u�?��'����͵_��'��eV�~:n����u������{���$�S��O�~3�����W�j���(A�D�!@$��LZW��PP�$�<���n5]s�k0��\���
��l8TC*�p#�	�֌VD2�z.5���������C�y��NX�5�j�$�:6�����0��XF��4��N�}����G�'w���Ǔ���8��}R�ADc����$�i�itOd�פ������L։u���V�	��U�]zM�Je[������U��V���7l��C��ُ)Z��4�� �%�M�n���;�8r��*	����u�QͰ���ѭ��g�扊�b�k��2�ρ�-e�nhQ���d�!�NyG��R��ͳY �R�����do�:�N���4x�hNgk��X0r��#N��|Ꙋ��(��� ��[O����x��J��G�,���DJ�R�S�}d]�8t��~ L6yIjw���7����"�����
�W ���!o�� �[V�knѡ�[3F����BN��A�E�=��{U�Z�F_K�i�~�������)�=J���	�z��6�zq9N�y�Hth��픻��V9�e�� �_j�_���
z��`��N�ݸW.�6L� Ӡ��*͢���s���+M�Rr�͗M�B"pHIkkY �UЬ��%!��/�WW��6�7Ρ�
5b�.8�
[Uj�6з6>$��vɲ+��dF~\� �6�O��&iaS��nng�^�_M@�An�-YA���8vjbs-�վ���lC��xoE��7�a�p�zȦ�:�����H�Kۇ� �d��S�%����|�f���x�����C����M��V�����'N�a���"�¶�i��Xv�$g���~VtiU��xe��^�=꬜8�f���珵�-g%0O9�h��?���?�2�[R�U�5Y(t��4�����
T���'���E��=�P:�M�y�<'�E���䙚�VC��+��[Ԑ��7�'t�Vm(suy���Z�X�Q|7O\�b@­�@�с���pv��	��B���1-8��h�2��[�e?�Z.l�Vh��6����g
1�G�]\�Zaz`��K��d���h�Ju|�Ҿ�G���/G�^F�ϫ�d�T	�	�(U���P<F7�;{~a��H/��dK {��$t�$�V��c ���gO���A��X�	�9�Z�X��sB+�}.ͺX��͑����
\a�i�V���U��^�N�����V�\I#{��� �J�5��'Y4yyPHr�Rt�s�譽*�sA�E�aU�-�2���Z�,����8��/=�,ޡc�c�1�)��K���܈k�A�ޤ����,���߾���| \�U��N��h�3���^�2O)Q��g�*���:y���[��~O�*�5��7�W94�26�^TmY���w�_�d�)"7>8'DAC)���\�]������p��>%>Aa�[�.پ,�p�ؔ��k���82��8����xB���5H���l�ۿ�76
�V4��sWT�����C�̟����g=6"A�F��# �8E������V��ֵ��N��?�S��ޱF��o@/�:�?Po��I���Fe����m �
ؔB���W��)<�������pM�TRR�yṔ��*	G��m��G��d=r,#:T�y���+L��#�V�+#�S�~��=em��;ĉ__&ޯKV#�'����x�F�vxZ�<��5]>V��PV��I �J�����?��3Z.Ztn4�~��ʎ�7Ha�\'��)�͎�x("��4"�3ޏ8'7\.��/m��	u�	޶q��+�t&�H�䀳3�nex��'~�9vb4�r0K}��0#M��6���i.�N]�R��h��Ϳ�`������أ�CϺ�N���T�)�#B4y�e�LB�g�B��!���k.�b���Z��y|��#����T8�H���䧋� y{�akb��XR�<j�DY�2J^�@:1WUj�Ma�1�2Nr�e���
+6b Q�l�G�M��h�!"�o�ߪO�
��,|��Cg�/#�W�{�R�L���� ����|(���I�
"S�m��}z��
�.z¯���{��{m�[�y|�@`��e��y�Q��V`m`�X�Xn�0�����n�j�C���^U~À�����]���IV�)d[��ڝ.A�Š�C�ż�ogV-�k�0^�j�Q|Q��i�6�.JŉI|0h-�KȎ߈��BO��M2�����:�	c7�T�DT�>�33�iгg)�CEl;���k,��}d��tN	< ��H����Zz7�՛�J�T��ha*�(*�K,�K��[��_��K�{nm+�4��h|Y�>����@�}���j�Fv�/3 D}�m���ﶗ�e}R�%������G�m?Y���z�ACPn`��L����8[���.�\/����^1�ľ����^?�~[96gL@�D���&�
&T�8��'k����?����=���l�:&���*k�v�,%p�_���F�J� '��aN�r�q�"X��i�7cB�9�) �, ��dki�eJ�ӌ��a��L�M"n��9��Mu_!������uU��RDg���>�(�{U3v�3�yp�e����6�o���z��:�����~�7�X$����Ը����<"�����v��a���
uݞ����o�v�qT�&��Է�1�]�ߒ�`�X��$`L�����1�o�j�U��#�	�`�,�R9�Ll,�������_�V���vL6����r�6�*=���,'_�Y3?��w�{�?�p䊙�BiH��I!P�&	�5����ۻ�2�r�����u�1� �P��BQ/_ﴅ��~��=)�X4f��kL�C��X.ඍv�ɜՈ�J��Z��Y��[�������\}`�M7
��e@�M��j�c�M�����G��4W��M�%�����-��n�&�ޜ,b"�@x��x�4�j��z�h'Ã�oh+ۈ>{~�̔� k�F���gasY�%~��BW��z}Wsֶ'[�~J��93��2K3���膌X�ٷ�f�6���a?e���#2��nt�ҿ=gT ���n-%���L�0���a	Vt
���:J$.t4�WSxs�]s�h� �ٓ���V�|���T�w�D�X��T� �B��|�S�����~5\�.j��/Q�s��ݦ��@_�������wɟ}`�78�,9?����L��.<��J4(bx_^�>L���I�:��o�v�+�oO��6lj�~>E>/'6~�����p���dT ���6�]��['�rh4�P���~R��A�Ɖ�.��!���ϻ~']|3`�7��k��Ё�/�7�=G'ʁ�?coa��h�Ve%}<�����l�o (�*E�5u�Es��@�▒|ʊJ��ֆ ��4	���d*d8%3��jBX!K W���9�o�@���X��<�R�Ԩ��'��[�"P+h�j���=�j���V�p
b��g�`cg�����M�2��l�y���9�e��������qv��(ElpU����f'�(< G�������Xc��g��K���/�vI|a�ekL���Wk�s�� �:�{3#�Z�$l���Ɠ�EB`Ć�搅��`�n��k[�H۠.G���J=�!�3L���c@�E��\Q���bL���Ewd¢�%/��v��� ����qi��c���M|���5фG!|�v�A��@^�:��X}��hE�i����Π�
U�U�ɑU�tɆ]�����X9cb=�{��f`��м��'�ĲO���gh��?_�vp�
�������L)��/�L�<�iiR.O���O�!�Û�3U_Y�jl ���j9Ak��g8iD�U�����*��sħ�z���s3���a^����#��1��u'��q!�{Ͼ�7��-=�/���s	%}�|���0,�=$]�g�����-�@?k����9J�w�%���o��6#+�2�G��uTr�SS�eVP��ϒ�Z����t�P��A�@t�#e���U|�R�u"@G�nk	�}��Y)z�I�#ɚH�c�!G3\fN��j���!��5��}����]���@)�By�<��vrZ5ū����V���"u0�-n�)�~���[��w�sj$�g�������S+I�L-/��� 뙁��CC��~�y�3snH5�3W�4^s��
7�ݫ�����,�e�L֗�a������h�}7m�w�
-���.�,�����g�k_<"1ǝ�y�`%A�j���s�MnU����Q&{�cG�:�����ӫ�m���O�H�����DҐ����5$��$�4�-�����?�Wk�͇��r��g����ӯ��s܆�wv[���v�OuH 3$�Z��S�z��i�b�ڲ�vu=[�=�=�`D�!�ζY�����(@�	w��,8��G�uU����p�B�>�7�I����ͦ���9R	��o�r�f��]é;k��8�|��9_<����)�wn���#Q�r�R�">x�%A�0���;�	����:�*�!��cP)�+�jiw��^�γ�5&Tv}~��dpE"��6�������%T�^F���+C�2��)���e��C]�HT�����E�8�	���F��Ѵ|uJ��rۋ�tYȏ�\ˮ�FfD���T�J>ibr��.6Qy��`M�����R�£ ���PP�H.�
n#�NN��G��j49�Rj�b.NޙV�D4c�+�2�s�@z����xZ�{>�̫<R���?��x�C�kI�V��.�s�<h�J��M�������'��_�X"������eD�GB�,((�x�߈ȈwG��S^�M�`|jz<��Ѽ�!��N>0������w�A�q�P�i�?
�J�i)eO���a�\�~�*{�c�q�*���-Y�ܛL���v-"�eD�mmq՚�ݷ�\PPժL��"�"�4��������ҭ���ْ�qoDSe�|��V��������)�`u�F��|�<VU�x��n)#��g��:9��.`��50�&����x"��=���x\��r��y�n�X*�C�ؽY��C���h>�A��29◍�s[H��t~�0ۇ�Z���v����$���mu�&\����zk��Zb��Lɱ��'d��8X܈�k&�l=�/����|�'�:�]㱵��ǚ���g
�%�R�OxH���~�u�Z��)?�L�sp���^�C��^�\�(B�cp���B�u��^�_�&��~�6�&N���8�v?LQ��"��/��
Q�S@N��H��?���Y��O1�-%�o��EI�̯|�N�!.m�g����Xh��L_��9�!h�()��䓎�~����=�̪�Yh�5��L6�9�')��hV趆�l�O�{�yW���"D�w�Dko���*8�Q���j	���SN�٢�b3�.�91�������!�,f�Z���x���^���t�+R����T�
 �2Q�~�@B��d��bd ����p�jCx�X��{O_��V����'�F��mX�4 �kR���3�K`�p��
����Ꭳ������*���=q�u�ٛ�b���q�摔��mG$N��;���u s�^��[��x���R�f$E?�M���� 7&��O�;Ǭ�A�V�X��T�_�Ai��2>-\�@O���K��@�?��fe�{ٯ�`�-(4fN�%E֏:϶V�4E�L��������<�KZY���;5V��%��#�d� �|&�Gx���p�~�w�k����sV�u!���e��+�c_�>ѓ�[F|��(u���zV���ѩS^\l�� 8��m{�u?�w�>����*Q�{�Zgo��^��i��=)�y|�|Z��e��Д�2di.�%{�%�B�s�B��U��?���R�ٔ޴�gz<��m�|C;c�����D:`���-�sb	n�n@I"Қ���@�~��2WA��3��A������6_$ �LD��%�x)��9_�ā�!�>䭔���l�+�%�Iu����k�W�	���)���2~�c@o}zk��7|�.>F3yE3���1�'!2�m�)-<%���hڷ����E�����gO��&�_b��vW���"۩��'�=Ӎ��~7�W��gMcw	���t5��?�0��%�b��j[�Z�����ņcQ�#�H�����x�o�I�9�A7}R�}����1���|��8�B�_�f��N7'|3N��q� ��`B��g�I_���Q�;�v}���f����iG�&���ᶸNL2H��˷�jOPW*N�@�av�mf?�|d[����w�G���><�s�o����x�&�Ix2}��/d>����@R�p���n�#��Pǖ��&`��48���qս�_b�bP�=����즥.|�����+�nZ#b������4b�R��pcl���Ԑ\[�l{�Q�K2�[wB��2��fY�x�PO����i�A~��cqy���ljg#�[��� u�-�=������K�ܹ�@J;D���L���� �R~H}�G!ι�Z�c���\\��|M��/�^�U2��ܶ���n�G!Ī�	)�
q]N���4���ysC�M��ZGV����0Ư�ո��c���(�yJ�w���aj�ك��cD%I��?�B��R�i�G<����� ���X��#�b��Aj�y��S!5˩���#����؋�q������c�Da-rm��Kz�
=k!}N(�Jc��]�#MpZ��2��e�b {���lAO�^�x"�l���g����9l$��E�LEDh�!�~TD�K�&�DU0{�G(��������*^�m�� }���u��[pYHeg:w�˷���V=D/��	t�Đ��64=l],��U������!����@dЊYa�sf|��GsnC��2I'k���p�e����J6���¬�-H3<F�e&?�`�݇ՙ{��O�cB,��;L�X�.��v>fY�˙�Z�pl�e5�E�L1�X�������Y�a�/	9^�(�����[Tg9ф�~��i(�e�����v�j[~s�V�`��@�3~��P�����h���I�m��W��w�7����wl�����G-b7�{햂4�m�������Lj�T��p�G.�j_ȭZ ݮQ�¹W���!�Ǖ���:y�1��똈G��M$BSt�ɶ1_�� w��FR�f�C#�EB2�q闾p�泒]�;��i�L֛Ϛ�v��3�],lȏ�S5o��v�k|��n�s�lޑ~�챚7�¡o3��1� ��
A�(���ș ��}F��;?���l�LD�16��)��s�D�Ya����X;��`g�ⶐ�/>}^3`�|]�I/Ü&�5l���n�϶�����.�"���v>u\Z���8��Iq#��6���k��_�:���gBS�I#w75e}�U�N�����U�6�� )��Wǯ?
}�[���ڇ
P���愾�Z�ܿ�:4VT��������Ke�R5iR/?�@N����w�f~�����=؈�S�WQ�ka��NGo��<��"�h/;��`Il��ޚNs^�p4����x�-��R2�N`m�}\�gA��]�/]ӌ�#�P./�=��y�8���>2�� k�#�i�_���Ll��.��f���Њ��yn/���l=�$�'��E���	]��y�BKI?29�sD��xo`0jAJ0
��Bz@3�QXD>�^�Y�(�8�sc�u�m�Rج�&�:Y��b�|�2G���� dH� � �[�u�KB�6d�&J� CN]������պڄ��;c��Q��с�u�Cy��o/��hoY�]q�.�R�U��e��P��yJ@���
�.�:ȡ�r-��TS�㕔ToU6�[�/`G�Q�CV!�\��W�*B��/n���9R��@�B�Qà�ރ>v�$j��Pc�R^ǄU��[�{ѷ�&�*B�;^V	��w��FSA�Wk�X]��R��1��Ȭ��畹;|���y
);�0!C2�W��1zg�jr����!�,ӓ�(MN��He�ٚ���f���[g����;��`���U0]'n�
��[� XPV"Z�#���ug��4�;��Yz6ax���t^0uqL笽��	\̴^�wbT���\D}�q�L˞g����
�M?����EJ��=����ӗn�6���L�Z�ippuD�G��I+�%�/����s���d���O��eR���7��G���Qa�{���H���	����1?X;H�Q��Jd�Iǵ�{�P���cד��,tfo"8���!rM�FO���ρ��6�^��y
��[��y�N��L
�����������z��_L�\�;�s�/M��p�hoC� @����/iω��ɶ�6�����~b�.B����+ێ 9:���BkU�����|�#���`S������dE�;�$w��7~�-��M��H�V����,�NhJ	����QS`�����=��[��@g%'�zJ%Ck	�9�.���2Œ��[=�R��1Yo����v=H-/lW�J��P� ��:�|��v�Esod��b�q�m�;�]�"`$w\�����>�?(��О��|S5��Wj��Yi'�[<t�(QK�Ͼ+�;ǟ�,Z����Nz��&~P&E��� �}~�"���J'm[D��J([i��F#'�Z�z�(6>&���&��zF��L��b�0�+�Xw���JO[�]��A��Ӈ�=<-�AN$�k���4V��T-�|�u1,�RT?���_]�q��/e��<ی{ ժp=^�.������o�M(�Y��c^�.*���0��ʦ�8���:�r1d� ������#����ɓ�0����}̣��,��&�u�����N��:l��E+y�PP�r���/��]����S��_oqi��j�i�b����L\�Y%�+70Bf��]��D��W#�?p�ә:�5��9;y�$B�� �/:2��!���!�ĮQ�ȱ� 2kÀ�l:Z�{��Q�V��=���^�-��P�8PB��6�K���ې���|�.#wz�$o!,Ae�N�ص�yO_���U+����oN����XX�����T�B��7(�Gmc�$ ���+�_v�?�gnm�%[j�>� �uwĉ�wf���&����߰��&�Yx�:�kw�(��%Y��hX�w�>]#�9u�?�Tg^}�]���R�I���RYN	��G;�<�>���Ƣ�f�Qk�ұ��[���3�n�u�e�figM:A#,,�Q��x��Q�=h�q[>ٸf&��	N�3�����������g8��n�O�&�,J�2<��e �q�O	�0Տ������͛�UG��Q���麄��?��<��`���=b���].�i�g�79y������/�q0�b^~����hvbg�����Ǹ�2����-��X�@b��5rSL5Vܳ�iG�2��n�-�g(A`+n�\\1����6�����f[`��Q���Ȭ�s��M��zu��5��h����~�')�/��\�\^f#롧�5�zIi��o�AE�� D����b�sz�8�D��4wK�:�jk���.�
�ζ���f��-�.\N�=�G�В��o�Á��?SL%��t2�އ��m��28�3�� u��b��Ue;׿`ɪj{]2��'�yNj�E���I��Ż_��=\������
=�h�.�Ù�9�ҟRE��'y�>	����4�C���d�2?IV�������|;TLX��4�Ä�����Z�'�Z�8I.E��� |���R)��;!7�������îp�f�6骝��pPR9�W�� �]_:D;����Ƴu��G� o 6�	��=W��ao�\���5>�oJP���r�mS丰l�7�q����l�m��x����=��Ϡ�6b��B�ܧ���:#��c2%G�<H|��=~���Dn3mPԀ����;K��J���X��oW��/N�\�<����lIG�[P'B�Ε�O�O��^.,fo*���~��(7;�F(e�2^��7�������6�(~������w�%{�"ŧT����U���� �1�b��Z�E1h�4�+��]�Ʌ�Դtzd��<W��'�� �`J�1%�:�db����1ўAzWrN�xvC&zPP#t��,�\��L!�Xf�:O6_��;T��}�%�U��y�C �u�r�"���Ɉ�U�&��Z �=��-�H~;�x��g�|@#�����ŁO���o��k�J�8x�yyx���g�nC���?q�p�d�8^��"��s
�Qϱm���8�
���2@K��~��J�r��:jH���q��gy�;,���ݚfgE6�6���k��^��5s���dj4�9Wg�� �#k���
�b���hcf6��R���mY ����:	��0��"?`bh;0u�9ިZ�� U>.�ܸ�c��$&�ϓ���u�U`��E/W��	�����79�����N=��ݫ��Q�b�����#��A)� ҟv�[���Z��.KEc����I���9h��
2�7�<���S�n����̤Gb���#.���}�$�X�eZ5+�#�̭*\�f����_�Eb�.�3B���NQ�/G.B<�����؇�E��بy�X�>�)8��r��]�^�\�!d����!br
e��^sH�&�y�sE3y{H?�u	�_�CFʙ3V��Иt���⃮�����y���eZ	Q�4$�V95��&��%V��oS�D�\!�m���b����ݺI�.��r$����+�hDo�4�Q�`�}���JƊ�_���De�@;��T�O�NO�{ �&��)R�}j��:�E��T���e-�&����ԯ����z.�{�$1�1q}^��=K� 0�i��DJ��^!���i�o�k�a��vT���V~�k����q?�,ˈ�崳羮U�0��S�¬d_��YTj��8�Γ;߶�
8M���T~t�Y�T���O.�^Jԫ�����&J{��G����M��E#��5�β��Wza"�:���3S�L�hΧ]����C�e ��t�^�\A~}�#0ya��ydK�L"�:�Y�fV�{���h�텲>��<�Ci�ȋ�U�G �'f,���F脻Թs��gp���2�J{ɡ�'c=�t�dPk�=:4X蔲��:R=[�������:����J�{��� 6�~�Sq�x;U���PݨM��I�h����m�����������FH�qA�6����
���=m� T�ɾ��A����Fx��^����_�JQ��	I ��w��Z3�{.�x58?a�K_��(g��ACn˘xA�ӡ��5n�pd�����9�E#�ΖN5�a0mN��?Sj��#���+�Ƴ�7�
���|)
m�~I�xEW1�؉�]O��T(��<�K��?u�jY���\��0*������d� ߸>�|E�����㩟������������}���[v0B�I�g�����m�F�B�,X�I�I�����)d��H�Q|���n&���Er#?�Bɓ�r���8�r�'fI�xaR EK��\��qju����>Y�_ڙ�gF�؟lk��������;Mi�$&`V_�;� 2Ԃ�w:��.lm�n�<Y�Ņ��C�d+yi����ۥ�d��=B|��(�5? Ƴ�/�f[�nuh#��E�R��ٽᰚ��^�	XE�H\	����VjūH���{����l����y�NA#�+�atnG� ,���Zd�}�!?��Gz:-d�q�Icpf��p��������~AE��g���D��oq.#׌ފ��[���`���%S�d������ �]4�Yp��
@%g�F�P�D����%��Z��3)�%�Gf�����DpC�C����JrퟻX� ���|����t0Ч���buN��<��Z%���y~��D�nu��.;_����7�$�E��)0f`���	�d���٣��U��Ȼ�xtaɬ�.��0�畬/�bk-�Ϩ��ںs�Nr47`���r����"j�.�g�,y%C��S�|1ۖ����"*��Q�qe����3.��5���K�O�=�]W�p��5s�g�M�u�)V.�Ԥ�?�2Q��)��/�nEC�
n;" �f�V�%E��0��'�<�T+d-Рjõo�EE�Z�6�
(#U�&�w�7'��*���b*�ob ��=���Od=-��():���)i��F##ޔ�2G����1j��������r,�r�N���M����r4l�]t�P��h�9ΐ2ж9�\�J5�TAh�_{+���$��$R%�"�y��H_����%I�A���������E�}����G����M#H	�d���hd݆�pU�%$P�)�4����w2T���`�ɟ���0��n��l��|�B_��������NJ$�������th��U�=��w�dU 7&�؀��9������jW՟��~��H��J3�(Y�0+<��ٗ��6 ��˼7p ���g������������������_^P]��7��:����G�j[|�d�l�TŊ���EZ��P��)rUiC�d��}k�C6ߞq�ED^=��g���������좷��Jeو��E͌~���u;��z�ِ�b<��]���"L���
���9f��_9��M�8e�����1�ȂP�_��}`���%M~$��V^ %'��#�X�cU�{SF�{qv�M��=Ǜ�+�] B�y��u-�Яr� �_��w�`g�Q1�l��t�-����RrY��ĭ`p�;����{��S{�y37ߵ��àɄ�]~<�;Z��k�}��,skӦ���G�&�4����d�)�9���bM���j�jݭX�������1�A���#�{���j'��r*�qd�=�]2e!��lb����4s�X����m^s��^�������w2��$�:(ܨbM��u�-l�3�LN;���]�-��H�����Ѭ�9���9�0�������jX֋>H}���C��h��ɸE�F~���R>JK��d��]��E�7[^����VfvI~\�fD_���}���h������-�&h���F��4� �jF��K��5? ������#� Z?�_A��f�bʴ��4����-�ؤD�j�g�ם�0�v�F���T��� �if[�����3�GcCT�MͬD0b����d���-���Z@��L��*��I�&���W�X��H��!6�����2�S����B?�$�ƣI�/)�V�@�/t�9]�ű��I��{�)I��	��s�����`6#�A���	�I�g��΢�$�(��Q)��ŉݥi�_bF����E9�up�b��΁g/��nf� ��e�6��*�1�^�h~@��Y�M�k�v�ki*��=��Ng����"]LNSg�!����b{,k���%�o]?*]q^:n��Ѣ�4�]ãY�-��b��e`��x�ڗ��W��ɤ��t��F�m��_Zcށ�Ŏ���^6�3�x<!{?!uX'.�	"1��.p)�L�p�s����������f����1�o�����,H^�_`��a}�nӫ޼1�c_��#���"w�|P����R�5��1�rN3�����'��r>	��'���/6ݝW�J%�n,UI�jѬ,
}��]i��w�t��:����>e�==cDXK�;�+���l`��s|�f���������6���<�L���'_C���ii����`3�uC��J-x" -�W)���*�c�����/N�~�p3�#d#l١��	/�4��8U��C��Y�&(=&��k�ˈ�(���a���U6v��]wm��t��� ̑�<� ��v���b*�%��d喱��[���g�[�)a>��˟�i;������X�� �u�`t�����yu[~��? ���0ONUb�;6Q���yJw}��_gX:zYƵH����
�������ė���y�Qύ��2ی�r���5�L�P�����û���:�V��/�S�c7�<�(,ϐ=����{j�#�����f$T��9���D��	K˴/܋���PJ"�`ױ���	��������}Q�p���HnT5��"3�h�s��͙��^-�����V"��{���7��v7k�@�/Y����)�� \���96^�gH;�S�%w.}s�^�vK�M�&ˎ{Xsu`;��7v���|*��se�8���+��X�m�6��/������i�'��T�ӱ���dj�,Arg��_U��T�w���.B������y�>�W��so�:]�Q�+9'���ǲ�~7rÉ�4v*���t>�}j3�W�(�F��=*� P�P���5�*�=�^���]�b	~PHn�p/�'F���']�V=�.X!����[�}�}��y�1�貥��0N���&Ư�Ю̑92H�t���#�L(����F\��Y��Y�N��Ma�:F' ��k.��3�s!��E�PdB��b��*�]=(К�VsE�Iw��ϕ��I�?�ZP�#5��`N�G�=���o���_�œX�	��0��\gW����v���S������r�|J2�R���ö+>���&;|-�r�3v�0W�鴠��B2٬"q���ot�r)��KFEn<���,��o��x�*��|�9f��B���i @�Tq���s�SA�3�~+%����e%l-Z��.~����E�Ty���(YS�Ռ���NQ��Aj&�<X^��ߨ��0�&?��)<M�����腶D�	?�&R��4��ޚN(��� ��j2����Mbޚ�3�vɈ���U���D��Y��9���2JD�۲��o����D�5���0��b8hi��3x���ذ!ކ�d�$���5C��?�;S��n8=ؓ�	��#^/*���p��#�:�~���=����|�7h]�.���Jgiՠx!/zjJ�b���JT^Ё�\�Ǧ��۾C[�	{�����e��\�:�@���S�[E���zpr���Q�;�8ö�m�t��P(V%jUZ�_ި]����g_Fj��oz��G<@D��z��`����D�
!�c4k�x�=��7x�?�]e��Z5�<4��Sb�d{�1����طM����ޠ�:m�xI���-�G�̻��$�|���3L�&�����͇I� �Q�@F��v!�J�$$D�&�0��f��Ůy�i9&'݊�9�zc�R�}'�Ws�D#��/zq�<��W��QL��N�����ޟ���s��<���m
�@��c	�����,���c�"2g�R(�:��6��|��ǻ9���<s8�E ߫Q��#�#�r���Tk,(9�x݄}i�_�-�������6h��
�&�ؘ��~1��X8����16/��Gq�wû,�Fs�+}���ە�\<Lwm���'3K������9���wG�ũ��(rb�Z�^bd�\�EY3*4�S��S���%;xg%�������5��M��M�V/�Pʃ��i��`�)�8�T>B�'�"��PN񎇠��)g��,	�>"�d?&��x��,7�Z����y����9�%l��7��yCΨi�_J�,8	�*�\{�@8�Z�;��
�c��w��C< J^���4�4�g�h~����s�S���x�Q��5[���{2aE+sÏM�5���=�)�iO�������!���-���vZ ��[����֕^��a2��N�i�+c�"(�3��J3L��Ib-T�����}�� sA�L
Kw�t� |n�hC�A� v����8�,P�K ��`��� �c��{b���ڹ��]�-�o��z������J^>�<�����..1ʸ����C�a����'���ҿ�ƅ�c0��[y`��Q*$N�6���7C�-
tùu�%��
��b��~��n=�����+� (�'�LU����ˠ���%Y�n�[�*@���DGb|���h;L4|?����|K$l,�d�
%<П�Rų�����)� �*mk����Mr/��!��}����n�4����"z��0�EDmRLL!=b vI�J���)B1w� �\@]�g��瘟pV��L7˿��U�����h�]�4��e�C3�]���ډ�la�(�Wk+5j�/�"���j���^Y�l��ܮ{7��4K���=vlr���������P��RB����U�oK�	Q3NY�����⊟��,4����olU1t;_�x[+��F�Q'���.�yyqYӽ�/�z��z���F�5���}ҿ����kzzB��E՘ʚo�đ��3�����qt�jCP�"E����2�W���Y�/�����B�������i{An�y$�_4�y�� s���2�8Vg��2��F�
��~h�ڜ���/�Q�F������ʔuۖ�Cpu�����6-u}�~���Pa��D���ܼb�N<+�E�$��ƴ�xݞ'��u�x�ͦ��,h��^^]�&tNa-�tG����0�x|��S^����5��bZN�[a��R���`��>\
��!��-��t�\�RN}��g�_c��(�6��^����I�iƟ�*��_�+�>~���mti绷=-�I��ՉӰ&�w���黬g�=J�Վ����p<70Y���&2|�����+HI���	h'{@�k���h���כ8�Sg0�����M��ѨPR�\R������\���_�52`��S�%�D��(��]
C G�m�OA�j=�`��?���B�o!d�"������}�{,� �0-��gD@*Πb�b"R��}�����f�@��i�P�
��%S���z�"��%��l�����t&<�����4���=g-�*������L%����G0��0�?�w*<����?����=��d����((H�W_"CQ�i*|K��_!&FTG�ч"
׵�"{�����C��&+����_b��KCu����hth�d��霥�[rѕT�ҝ՜��]�
[؀�[\��BT3�(65�٣ )���PT��
�^J�����[�]3�3@K ���?�hk]Ll�ݹ	�<FrY�vR�>A��2��e����i���QIc0Q!:��݁Cdi�_`Zם,�H�W��B@W/W�;�w�8=-^ݦ��5�z���l.�a̬EJW�72ӹ��d\�6�����Pp/�ꂬ/mw�(��f<�7��U��=��uT�����������m��G^�����	p!	׭+����3C�K�QUC��лы��Q�b����y��s5���^(϶0Es,��"��φ�u3cP<�X���v{C�����u��dS�"@*�U�P%�O���W���X"��x��O�b�jQ��&mda�%��{Ĺw@J�v��g͢��Lv$��2k�E�@�A�@����V��R�^,�����+�+"cy�^j6pՁ7��C�	F���a	��l�w�5h��Qݣ"w������z�iٔ�ص�M#J� @���Z�����shX7��=j	�.$G�r�>�$�� ȟ՛]�A�}�<JR��q�*���K��G��k�I��!�|��3��/��k#`��3*ǚ�>��@�CbVy[��1Q�����Ih��HR�.��\�MZ�^�_T�j���%N)F�̛Ä:)�0;p��� F������&xgS�h��`��ju����ˬ힝�q�Ub?ٶ�s6Ӆ(�E4��Y�97Î����t����Z_��|;�wD����mb��U0V�փg��Ò���$�+�sW� L~�`m�m��tX!�(��um[T��w�Q�.@�gf���`7�?���^"�
=]2?V\����!O]蔬Y	�r�z !7�d=Q֏r5 W]�V��'�=[A�X3�CQ�@;��C2��xK�U�&|9�Ь��.���l&�ECP{K%������񊭫��\�x�7���FL�J�6�|�*��J��e�����CH �n$r.,'!M��q�I�~Ut�H^���}�bo�o�S�����,��ԙ���co�a�qV�kx�r�?2K;О�_kn���o�编@�43Yؘ����sp3J󥩬;���R�*x��] wp��8l�҇�\!ӷ�\,�G�i�&�`���^�ȩb�Ç麾;�������ĚSc�Ϣ�(k]@��(�X���sh��:?��RcoX�l ߦ�5h������C�)�(f��B�@R
DFjQ[kٮja�}$���ޅ�TVv�oP�I��pt��Z4��\ԍF�H�6k�^;�������(�n3�0�����m�y]����� zq�fi���HxΡ?/��pPS�!f��_���ٽ����j9`
�~1�zf�3�<���QUd�ɖv����6�yrk�������-\I�ؓ���p�e�����B������+����������2�
�*�-pN��\;�C3�-�+��
���c`&�;�X֒~�6+5E�R�ccl��Oc�=�-;�ἅ���j_j��C	%B��׻�Le5�/��_#{�!�%&��SR�1�L0*+���9\c��	�
���O�����J�bNn����|���k�9��skoT��U��$I|��Epc(	ABzh^.��U���q#�#%��K5�˗b8��*�X�3�\w���7���!��ŕ$��|ƥ��k��f^7������oR��1�44�3/�D�F�	uRր:!_('��[U�1��2�6y��$����V����Y8`��3ze.��Ge���yg[�@}W�rZ������r��N[I��T����vq+F��r�˺���|ۿ��]�`�z\��i.<�֘i��Dܵ�4618�SyP��tLa����5T8t%�|t}��A���H�Ʀ[ϭ5����=��!�V/�g�#�ۿf�$ǹ��d��0��%��o��!P�,�|(���k:�H%����@`0�-�ZoR�����G�K��vݸZV���ŨU�X<CB#[������ ���@�[F�%0N�
�]����gG�}���5�Q��s�`�|@5�]�6������B�r�{R�Yp�zt��By�cts��]�o,���=qƦDMsv�:��#O�ӛ�"��"cr�2�o����zŘ+E)�5FFHkN^�����e<�ŵ����2�]1�߆�<QcǡP4s��PÉ��4�{��-�P൞�"�>7�]�"���"�61�LD���~�Y���l����u@���%{j����+��l��xjtKD ����\�H�e�鐝S�y2z	w�ѳML�E1��	>!�.���4X8��]i�t	���o<|�O^t���-ne��nBg�4}��Ć=(= j�p+��;P��3R�P��ҳ
��b�c��q��i"hYvnJ�W�*o�pg3@��g���׆
#�2�ÌtZ��b�hPE����Hz�7�S*�I�2�g{ԝ��W�Ñ>-��&藭l�{��[����.3�]�u�ʔ��I����b�n�3Gb�k4����X_'N��-\�5��@{QC��C��3X���w)fa%��[���"JhH��4�R^t�:_M5A��NtĨ��)�,�ޢt����|�*R�U�3�;���Ybv�������i௷�2��Xn��:��c�\�^�ZU�y}�7xE�"�u��}dݘ�"�]�:*+�S�A������}K;��x��;2���*?8@���A�o��� <=�Jo���V��)#h}��s����e�(��⋟��c�3CP�i��|���:V���6�s�*ra�@w���6�4�$R|G��_�s۠}Tu,RKV}	��^$I"��$�,�V�n�����f����� ��-t�� ��`K�^, �G��թ�ez�3��_�`K�_��
�����\u{��6Æ	?�Z��_kWg�!�����*��x�般�x���)�����s`o�����4X͆`�3��8��R�S���<�O��g~�2�j������_;�b�PX���v6@@�V_ɢVG�YW7�	.��6V�OE�a���%�r7wd���h8h�1[�U����D ��ӻj8�4�1o�pH�[/G��4�K�ݻ4�,�D�x��U"�G?�㜗h��j�]�# f?�j�2N�p?�J�����7��FH��T�cL��].�6�[	ЌLy�>������wxi����,T��z=Hj�/=��T���޳�C)K�0�4P-�3hw**x����B�����	�dZ<���{ƥ�B�8�/o�mJ�m�Xu��4
�E"R�͚��Q��N���Sȗ�"�/B��( �ә�p���hA�2O��{R/3����k��S�+��6c�:�Ƅ�힆�G�ښ���<��dc+
�	K
{�;�A�ب;˦����%�M�ۆd���+�A'�H.z�!�1z2������	ߡ��E������8 _��QK~�߭M��#1�P�O9��7���n!�>��xò`X_@Z\BC#J{m��~k��1aĂu^4wєC�L��L�籜r�o���SG�7���p�+����Uȯo��E˘�TgY�^����+���0e���P�{�9ج������j�v�:}����SWa����-fK��]�=����K`���>�u�j��p$�e:���r@�/��,��^��#��ޮ{��s�ii��sbX�^`S>ʚ����\��]V o�򫸣�!o.~A�H�5
�Br�Mp`�G����X�l��_\p�EmX-uY��Jҩ�<����Ը��h���8�fX�?�Z��c�� �&q���p���! ���Ip;�_+�^���M�ٗ�*�q�89���3���)������Q��s[��7zF������&wWʮ�5ٻ8h���Z6	�����_�O�����#5����kyRn"�Zh\�.z�e@���"Ȩ��slswz@o$��;��=��3�+&a 筣98�k8Uyb]+�?�p�N�}ϵm�2���z��i���#�--@d��yR�lN#�&�+�G��@٪Y�S�K��M�@��&���G<;C)�b�_O<s��5x	�>������� �
��U�C�>Za�4�Hj;� �x���o�u|Y;g6�0W�-Tbf4��\�ZY�g�9uE�|�4u�e�tȀ�t�b�ctd���"
~���h*k�`�P��zG���b<���΄q�R�fg�R�S�E��-1>_zH���O+P�}���� �����ƴkƼ�*6,�qb�ɡ�'���
[�!�=���-���̼�7-e�k���1�7w�QEW�.T���N�?5��8@�.����y�s_R�H�MC�G�#H�g=��Ҍ�<#�����HM:��ߌ��O)�+��P)99V���P !��:���1�;�gzs�kwIj��6����>Ԕxƅ�\U�U
��k����0���ܫ��Д�j�ֺ��x�Ȫ��r������.ܶ
������|02l3/�$tG;bX�jr��G_Š��kR�^�u��Z��dм�7��e4mG��.u�<�"�M��JQ�	M�]��h��' �o_���}��&m�DּLr>���3�${QB��O/0���Z���}϶�|̉B�ع��58`
�$�~���>���V:H��-t�K��ຂc�t��W,��y��E�o�S� �o�}|?�U�X�-�Q���Ȯ��6G�;@���v���<ߚ���%#	|�qO��P��b]9T���oM2l���F��f(tsˇ��c�P� 3ܣ �uF��2$��$sq��H�P�PU/h���5�3]+��3��~�>�����]��p�\�- �wp�[�9/+A8�^��pT�ܽ]uѤk���L)\<��V��$� l��R�P�U�Aj�������.X�/��u�7P]���_��l��f�h^�.ɠ'���nq��4\i%��o�r4 r�b���j�B�e��P4Q~sK�\�l��t��3?�cL�ӄεa|���e���9�5�@tg��i��j�+��A��y�x�x���q�8ŋ ٥�$�)G��I\�=܎-������ԠTY�(ʂ����oW��K?:�s����o��7�ۡE�k���f�����Ö�k�$����̯����@����rj�}��P��ɧ.��#y�:7 .��xtT��<2�M�W<3�e���*%�M�Iث�f��,��Řa�c�nH�]���>'N��~j���å�4Z� ��6h�C[?�& ~h>�S#!�7�s��K�,�}?e\��5�s��7k鮀k�1jNF��Ӄ%��~�u ���0�w�<_��/=6�2O��%#n�^g���5?��hwS��9�Ϲ�
�Y#RR�=���uM\W�,tM��	��J�ܙsW%6����B
{�Z��_6l�qz%r)LAT�@���͙�4r���J�e����ZA�c�`.MJ&,y����'а��2G`@�s�t��o�*:�Ld.��F�4H� �����z���8o��/�Ub���cz@��=4{:M�+!��`z(���"��Qq��Ù�� q!1bZ���Bf.<-��S��:;5}۸��2x�eXު.` �Q[An�<��:g��s-#�s:���(��{xI�e&�'=��qȠY�F(�Ҁ�s<bٕA:�Q\�_/,���N�13���M��x���7�X^*��Κ����`������� JC��nnu1���R��n�E����j��=��;,>�Б��s�1oP]㕙��A��&��)^T_V,-"C��a,RG���������*A� �@�)�6�飚]�Ϸp���O�.C_����٭^�m2Q�I��[�"���hb�KrGPؒEf��ҳ�q�L�������$��PC��W}��ĺ��1�W���0��\	N4�����p�#"�!�w�6��Y�زW�������/���	uU��I^,3�`�+��փ���,<n9J��$qсl�BB�,'Z���Ӑ��\�\1bz����G~]�і�?���{��+xW8{"��1n���@��]YT�{2��ر�4��e��)�B#@�r_'!{�Mмy c;>ϑ|�,O')�R�>x�Ci����]���a��Q�ݙM}�3� XP�j�P��2IG�>���҂��M�����m_�d�ک�E}�a�p��ě�m��ob��ʗ��=&6�kt�,Bŝ�ť���������m��'f��İ� Ǻ:�!�6�������	����Y����H#�Ml1
�a��:�������5��Ƽ�Q���:��{ ��]I�(�|�6�H��A2�v��i�`1�6�'�(e5zH�������h�[�N���4�OQT����^^a�A��԰JhF&�GeH�,���q�dt�M��r� �lf4�ʉ�bl
��5e���3n�mO�L�]�,(d��#�F.�%M�o�����w\��D 7ާaХ��@����@���]�����4n�BQ8�������yShn�l��ߪ<����(oϔn=1�㪠��q�2�;ѯ(���f5�ʼP�S��kɫ�1���ZOJE$��h�Iӏ�UP��3x�S�ԧMi���7�5��:%m����A�
-ȓX�-d�Ձ��>��!��j�q��
6����\	D&��~�`��h�1R(5n�!�+j�o����N�L��\�\�ާ�@j���HL»ǉֿ�ݵ��B�b���	x��be� J`�(�%��3@�7�ֈc��p7Uz��	9��I��L�=��'�b��[v�{>6�M�7O�npk`��c?��Ճ���2r���h^��ȗ�@�^_��c�����=U��Q��x�B\���*��F��e���,Y�F�p�fę��ypl�܁M�_�Z6Dy��So�-z�F^�Wܵ���b\�*�p����B�n���?�Wl�b/�[Nw����c�5�MgOՏ�p�meƀ։g���$W[0���ੈ���J����>D�\�G&4�kn�ht���a���i9�6�N8�6}�򑪮T���U"��7S腻A���E�aƗ��96��zu)U[$%��:5'��'�� s��E�.����}G`���x��>B1-����e����5(�o����S��j��r�jN$�ͻ�}��.���*�i�¼;c%M?���&y(!�S�Vk�W��mx��Pt��2D�O�D&��s�}"�@��n��̪����b��FJ!\d��^�ƶ�\ ����{�xGS1��*Щ�Cq?��&�E%���Eā�ڝ�]J��p5�0�#���Y���rN�b0����7��È��ƃW�P��3��t�T3��������U��W\:��+ո>J��Kmˮg(��w ��1�Xٛ�"8i ��R�vìu�<�3cW>|Kjl���BQ)��:?➟�g�hx�C��ه�e�ʄD�um"��C�:BNZ����2�NG�<l�D0>��;ѣ�O�t]> w�􍸗	/��e�ᎋ���s�271b�AD���ͫ1�]i�A�4�&�����T
vS��J�c��@�&�ND08�Pkk�|g�=md��(���j^��q�;r9�p��L.'d�F؎*���z�q̉��l���8��[c����Q�I?_�C�}�+�!�S��U�6m���Y�/������`W8M���x��(8%J�I������w��w�!R8SG(�����������1��X5ng�V�@V���/YU{�X-(��o���q8e?���l\+���Nތ%Ҡ?[���_}��d
���?�`�]�V��z�-q #3��WH�Z�s]7Oܙ��T����I��13��^7fΓ��H저�}�9N|�W3>[�}l~v����T��  �g�G������`7}�f��S�. ��%`�"�#S*��ӹ�;|�f��.���]g�$��O��z�q᳄R��� v�S�E���udo���G�q~:����ѷ��6 BQ,��"�̏���i6u0a���Q��ִ�5���X��M�����fo��ԜE�۶~bGPB4͠�����	�'�u-Q�".B��6���p��a�v�m?��c�~��j
�/�El�=��,�q���ަ���@�����AH0�>*S�j��H�qd:nR�E�fމ;FU疞�ץ��8��Kq�e�S��w�/��. ���Uˎ��~nEl��M-!x|`���V��s{i�:{��k�m��7���؉N��L���r{Y�#K��ķ�)\+�pi�xy�B2@����M�wz���׷vl�2�> ��@�ֈ���XR�r���,�y�A8�WT���?&� �$����L��pFƇ���9"��ˈy�O:�_��[�/� \���˔���������/�(P��ͼUS=E� �c�g�\>��'��&����_���$�ǘ09�5�L���7��>U���K^���ÊI���.=��Nz#�^��5�W\)�Ԩ�\�>�E@���[��7c���3�xWZڒW���H��x��
�aؤL�51A�Y�]�Q�a���� `(�5\���X��ڬ���'z���c���|�ޘ_�߻�_i;��l�tB���K�WNq7�U��ZD����y
�2G[u�:�����8�����9�8�: l[)31mVר-�V�fa9e@x�V���A�� �\%l>nQRN"_���0�oc�D�%0�ZeFh·l0��ij�h�B��58��Ǉ��2pTg��ѵ}?;�	���!�PR��C�KX롿�i&�g��W �>����C��̵��Φ�7�L��9�ݯ�ƭi.y����oX ��Xپ�*��p�ۅ���1}���)v���#0�o�:F�|6��;�>�cAf�ӷ�?0����Y�B�=0�r���R�U��W���Rh/���jخ��sZ�/��ZsΠ���cC�ebz7�\�@�N�m ��e�~?F�Ǭ�%���9ʧ�[�eˬ ���g]�qI~���f�Sa�2Ĵ8��m�ti�
�5B�J�;U�z%��s�QlL@��r����ê)��m�A\���qb��ON4���|aRWq3e�]��^�9$��|��-䋤/r�t��/o�j��_���HN�D^Ms#q/��Ƶ�9��w��}O_t�x9ԙ��`�7�C8��^��Z�v�R�T���D��˵�h�:ɦ���&�`��` p�$(��o��t`�O�5���z{��m˹�Af�=K<yސ�ϔ!��ٯKT���VH�}L��>��ŗ��e:djS꠸�����V�'#��'ZEߚh8�{?�:��w�:3����o3@�����K�N�G-)x�������l�p�C-k������[���M�>/
(z��������zw�����;����#������߱z�3����������]cٖ����@�̻(I0����f9�=���Sa($�L,qy<[j��_m���~+e#W�&e��0Ax8`�Z��1�Mʮ�}r�xĨx��P2�Rڥ�H����o��;�B;A���ZYBGQ�D��dT�}"�������Rb«�tH��t+݄�P���1bA��Zf+�4l�C����^�t�RSƒj����?��߿�&d�5�h��:��Ж�n����{*�r@���mՒ����&n���w���p�(���)�-��ܵ��w�e1)Qydmá;���C�c��:5���b��ęMI�s�5��OH��co��qu]i��b^�v�*�� W�N��p��e�I�Y�^wo���#�t�TF��ee4�m�I"�XJ�B�C]o}h���\�*�����r�N�k���}c7[����D��`�G?����	�m�\A$1�P�RO=mX�ꅇ��6�e avO�G����h�������֠�y~OK+Lc'Qj^XlxVHYEB    fa00    6ce0�.��F�6��ޠ�X�&����r���a�>�6,�&����+��l[L�=QQ�s���`�l�-r"4+<��<,��I�����E�*[%��H�"s�}9D�j#S)z<N�J�x�П�O�~�Z;�4��f�E_������́���Hk�ݬ�`�Y$�@HV���|2K~�/尔W���R9q<}Fo�V�:��WA��r�Q��w'�B2�3���5�BCӤPL����6֍&��&&��FM�0�gܒ�<�g뮂�p�MQj��'Q�ن�k*����5�֡N&�q��]7,�@�$��^B�G��
T�pa��� $~����Ջ}�yHR0�]Rm�V\�*so���Hc����CGZ�gys_5t	*��NL�,i�5�6;*��&�!r����~��Z&"�є�%�ףE�W�Ӿ������q0�e�q3���/�e�wU������"��"���<�ߜ,���=k��X�F��!�8j�uS�=�Ff��g����@�t2�Ͱ��.�1�k��tD���>�7�����C89j)|����ǈ�Fg�1��)����%��68��^?�_��#��/���9��8����N��/�hn��� Z��==�)G~t�k5��rF��az+=$eVx�W?���eB�Vzh�',�ԇ�Y��;��&~=ӓ}��Q%;�C� �G��(M����f�BԒ�D�N�^6�ʆ3����.j�3�;���?�:L��)8�d�v�R��f�V�9�X.�D�N��4��J��r8�jD	��Xh`��=ԍ.՗$��}-�X��ׁڧ����H֛<�ݗ��|6ݕrC��x�u�p?[u�h�i��:�x;+��}`dS�������wt�J����p����z�uq��r{!P�|�KJ�v���3V�YU����9�P� �.;��5g����bn%1[����	4Eܰ�C���]���}̋��wo��QH�`݉k��<�^Ɲ�
ơ/��d��ݮ��T�}:ៅI�%\U���(}f��F5��$�Ya�-�N�cn���MZG��-���^}[A����z"��;|������<�@Ef�k�)�p�!d�"� Ҭ���-�lQ�Kdqy!�h�F�\\�,WX�y��-H�s���vͶ����j�B��V��+�m�pG�ī��c���0k73��(µ%A�������g4`i�#N(�G�N�M��(�BIn�>%����#=�@�<�H�����ӽ6�[��BL���+���ҤjV.��*�Oc,��ƆcC�h�{������k�f��;b]G���j���;<�$��l��H)�\�
B3p�n�Ќ����e�� *ϻ��S%�R����Z~��]��Q�u�-U�Mj~gx�u�d��NZ���=�
��d�������;�(�R��
���%�[�\%hԈ���gK�f��Ez>(�{�M�B^��=�\��浹�po1��:�{�����Rs3�y�^���/p�&r���P��,fB)<�=�@�t?��'��8�z�tG���\���]6�צ�B��������*w)Po?Y�Hʍ`��Y(���w��� �x�T����.N��=ɶJa��K��f�Ñ{��5�ز%�����0�ZNn8�#mR��;����n&<�wEA�g6��im��Q��~�l��񇇗�ܶa���qɸv��ie��
�~��V�)�FC�P|����~��3���iM�����N��R�
���Q+��������!g���]������w���Ut�>��P�
����'a/��=�j�F���pϫ�Kx��]Q�6p�F%�-�m�4"�7Br�vRwR��캦q��լ�O��,/�`�z�d�#L�����8�ۇ1N�)5�=�j�JL8$N��� 5�aA��$���<��܊�����YT]���W��m��XֹW&�~�D9Q����QyTD��v�`��f��j��R��((�����
ET޺Z<��q_��)�I�Y��@�y3H)[I�[Uc(�0��Y�6��	R>k�ߘ���:Rn)U�#w���	�MK�z�U�
<��z��B�o�#��;�2H�m���m���;�?1'�E������l7�(������n~�b�Ac�K���B���]uo.T��5��te�subKv3*�򷝦���5ݓ��Y��>�ݛU��aUF^��g�׵th�W��3�g�v�ZfL�&��q���v�fcK�S��xk-ĭ%�D�\���]���/������@�$��,��jh$���m��6B�F0��,��-Թ�p.%�j�����9͝3{�m������k���/@�ESz��@��u47��Ą�j��PܐG8�?�/�w����Fl[Ո:i�"�B�� ��8h�hOZ�=W���3����sЛN8�*�w�e��JU���rd�U4R}����JԽ������0�C��hg�#��b:6���=V�����[ۓ�@�1�?���;�W[�aj�DQ$���R�~�`!�~�zR,|��?5��agߠDZ���0���!@O��Y�4D[�=�r�8)r�k�OŇ�;��C#��0�L�����>�H�:�ˬ���?��3�y/G�a�S�FSJ��@鲢�E�܉�c䴳ǟS��[D !>
�vV��ޭ��򶑱���^�F�����d�#���\�6  �� aQD\�^�h�8�|���
��8�̫R�5(�閞�K�G��[��~�R��H%.⌯�T�<ZU���f:ݏ�u��%0��8�z�qo��?7�u9�Iqu�/Qd�Y��i���	F���e��#��N���?ď8��yry�ѝ �a�oȂF�����]U5)��r�/��j�J%iL���h�s	�M0
aī2��(b��x[��L�?���q[��L`��߁����B����мJB�n�s��v�I�|b}f��4͑?�zh���{�������0����ӌ��y��8�'�V	��!-��-�V�u+?W"���_i�K��/0�ױ|W���#�q�m�筢��o�[. wqJ#TI9���l'�v�p�����%�ڱ1T ���Y�\QC7B;��ydSw�����	}���yբ���@�c,��W���S���
�*nf�܎�gOZ�^^����H��7N����;��y���Og��Y��J��������vN(2샍����Z�g��4K�$�]�&��:���)O'ZfD�L+�7��$��#�x�F�h-�;A�0-�a�wev��W��O�aF=�H��l�� 06,n�4��'v�	�ܢJG�M�;,�ѥ�rC��bJ
��r1��v��p �*�^^�������t�Q������|���MF�����]�P��e�.��c�+�yUM9��R@�n7U�hqr�7��"-���C�bP�����$�wiKu������h�\L��U��ڊ���x�u���y��8=�#W��I.U:!ow�e!`+0'�C�C�e]����ۢ	�g�r�2Z����;8���a+0^2.����Uw�0����3�īw}?�� �����ܝ��Hs���4�s���Fn>?��z%
�[a��oS���cb��gTw҅v��B�,��o2�5.6��#[)E��T���ۻ�����X����ܵG���Wy�B�Kq�n�#����㴡�G�r��wj�r9���-̣����7)K>�=��mͳ��'�x�o���;��5���cnj�iwl�*���ؗٯ�����!�A��b�f�W�`m��B<��pQ _�4|rܱ�Z��EG�L����h+|q�k�*Ř�	���i�&pXJ�/�=�K���}�OUb�Ҝ�o`���ڐ���e��a#)/K��9{�@�����;�!�'So��&�b�S%��j�>Wf,n�u��<H�`���Y�0`�m�Xz@�7�4Q�H@�Ւ��bi�6�q��1<.s��b�T3	��3R�C'��x���)�q3�����oZ[Md�E�L�z�fÒOFU�e�ֻh66L&���F�Wyc�I���O!�Lܔ��H�S\mx��E��W�;m��"�3���"��NF�p ⷧ���e��Nܗe�/7g���fQ+�j�����G���s�?���i$��X��B�(b�r�2N9��4�ܕ�:D�Cgk�2�K�Lk"�8���y���Auն��>�6f��� ��M����  wR�8:$�)�A/�E�����j=c�� <�k��I"\ �;��x��"��| ����4���ɵf�#��G�}y��J_	'�л��o�3�ٓ^>�-֤�8�/��z�g����N�cM�oB�?�fwS��D�ڞթ��u�r�d�b�p�W[I�4hV2�V<�I���أ��NSp�V�uz��|�cD��Y�H7�D`�J�|�{�-F�!
������Ѝ�cf��lE�����fe��F�����\A��Ȭ��!�5��D��H��c�_*�V)N.���X�}X����+�]�UH�De�n��BT��z*��� �}�S�3<��q� 1K;u���~��z�*W/��{�T��B�v�S�"%q �<U�#p�N_��=
���pp}u$,�H�%�P;��h�1�y!S�Zi+���-M�RR�q�6�<�Z��O���$ߞ� YxŢ$����zQ�'�0Id
��ӷ��fHD[�Cק�?����6��A �#��y��@�Zy�#�.J_�w�X�q�]<����w10Z����?,�z���Wf���a*���{M���7�K��[�y9��3����Fvu�ƽ���h6\��/q͐T�"��$�d�1��"K���7�i���	,�ڴlӕ��� |�jv[���>�*�ޖ�Ifr=1��J�j��y�'�:��
.���C�0R�(xw 
UR`� �s�;��Q\��ڕa�x_�GNb�_�L��F�<��q���{=˭m��WC�0F"[�@�#]ʴli��P���Ҿo��o925
R*V'y��s��Q�B�l&ࡄ2p���=�@��k�i�2륉�D#�|��!6 ��L�',�hg���-�>`9œ�\�����V������Z$rvi�r8@�����Oٛ���Ο������_@&�����vL�q�4yk��K��}S������g�J(�!��&�ne	`Thԧ3v��\ys�2V��	x}b#O�\�
�`��|�ؓ3�\��p�1�#����s�5�=7H��P#R���D���R���s�;�� Ε+�v�ݷ������DϬ͎��,�%,8�� {����a�������p��1�xg��4szӜ�p����V!h�d��\�n飠�
�/=Di2d�+�������B�hl��Z����(DOϡ�/��?�~0����>J��.����l,}v�ΊՑ]{؜��^��i!��K|���G�3(��4���w�Ƚ;X�#6Y��+5�o�dlǫk~-�O!�+��𤔤,z�*#�)�.8� ��hHy����e�>$�����"-H�aI5�=� ��2�l�'�0!��\�RV�0�����6	�z�5-��*�S~-�� :��Yp��v��V:62�6��y2>s�򶲒�@#�8-k��0:��s2������!6�F͓��-� �^?��2�I��Xi�P����;���r��+�ޏY7nUV���7ne��,�t֓.ꗻC�N!�fH��I�)�-�� ����x�� ��oaRl���%3Hh䒤@;�	Yr� [�M$�H�$���ň�r Գc���>ģH�^�t����M"gg�׹�Yy��~V��!*Kw%"�S��j�ǽ�(���5�����c�f�7�B�yQyw�s�b��񸯝䩊��k.m�l���`�7ң�L��e\X�N��!*m�{�z���L�-ӽ�����*ޚ���6��75��{���p�ʺ��K�i_�ށz1i�[#���P%/�%/e��ߜ�M9��f��~A����[�zta��<C�r�뵽*�N��d�f9ŤV;K�9aY��/3Թ�t��0��lF���U��<��T�t �wj,!��Fu�����Ƅ��}�zQ}�X}�DV&��06����u�m�U۝��Yu�\#�_���Yx��Z�?k/w�l ̠� o���w��k4o�_�Ht+-�r|줘�,!F����9�d�]���f\�Sk�iY�
�V�Zv��$o��4ԗ��5"��*W�Bf����T;!�j�s�a����f�@�6�����1俈2St �H�ML����sF�+y�7;}F�Ol��F����e��NA��T� ���CB�@�'~i�kZvt���+��f��bR%�;J,��K�ΘmƟ�B>�T�1S�iK����g�̣+9����/�X��A��w!a݀�x��Q��o8��DTU�=�����-�;�\e*]����c�ғ&�g�(���K��������;�HX��٧,X�PD�a�V-��n����"�`0� �񯸥�LF0:���:�b�Q�\t������!-���\ NR2d���L�g��*��i̢t��T���f�|l!��h�/a�z����%˿����b0:"Eϓ�f�&9Ɇ ��\��y9~j�&^,�y����_���oT#Gl��l>�D������M���J��� >����;ӍPD3�Jw�I�
�!hl#�,&ޚ�� �:N���x$����o8��h�⢕P��͝�xl)~�K��#�����i֙�2H{`Op�ߞ	���D�͂/�5���&2e����򥂰"�k}%.�Zr5�-ji�cO�H0C�|ۑmYT�O���=m�)!�����hT�2-1!��z�X�Wg�ͨ��Р�;��*,���p��졑 lB]޻�nKj���"æ��PG4�,��cU	��3\���WǙ3����H�	L�5,��4Ӈ7{Y�8�]C�7A�s��L�m	rJ�KG��ɻH�#q��焬�v���a�z=*n�Qn�(� &�n�[ �����5�%e��ӓ�6fga�p[9����!�(o8N;5�2�6��R���Η�bL���]è�y.B�f��G,�;SѬ�e�[���"�&pm%�wcʯ��3��e�D �N��(��\�k�����<��W�=�����p�d���3T�oٕK�HW2hi�n	t5��'9>����H�,/?�<M�pF��mG�α6�U3YJ����[5�nV6K��}��i���J~h��lv��C�H��͝���iz��a`����l#mޕ��(9ð+���0~��5�G����	F�}���O!�.k��Z��磙��>mI�vt��k�:�*��{m��_��D^�æջ��#i+�<~��1��#��?&6t�a= �& ���|�|,F@�������v�T����G�䶣��;i��ܶ`	����!����S�z��D��.���Y�h��ٗo�(_u�#�N1�c#Þ_� =��c��c�����ԍ\�"�z���}��|��5VU5ܠ5�2EDeU!dX���0�0��Υ��4j�%�J���G���Y�A�,!�v`́,�뒕�H�2is�j����������m_nh�2�p����t�&n@"VRu�*�v�%g#��*:�/ˮ�z]���Y�e��s���.�L�znZ(I*�辏�!���}�,sZ�L��f�FRts��I0�ۇ�w^�&q��o{?�'P�*�.l3V���wJW����IY���s��E���<]I;4r�^�*��l������z��>�O%K d1���;֞�q\
���6aTI��c�$FG
㿿�����i�Lk T'�7��qӧ��$����>C*�:��W�(��d��
.��1�L�%ҙ/�)��fZ�{�k2+��o@JWJ~�A�WA�	����?�`8;�+�f�����m��@$x�\�)65e_EC>�+������ձ)v�r�V(���Bef�:�x�5l_�/����p��!1,^;�3sJR�eK�7��*�_�����13,@���tuX�f�)?)��"nx�Ҩ6�m��e��xɋ��1*w>�A����&�+�og��:MK�]AM(V�zfV�R'�y<��]��,�2�k˄��mР���8��-j��C�o���.�+/�/���^O� ���l�2�qg�ɐ��y�xb� ���[�}i&-'�[��#%X��'��RHߓ ފ�C3�F��f�����H�!C��������<� ��qK��*trq��]f�(,�R�l�Q<d�HL��*�rь#�1�(���	Z�<����0���Ρx|�YE浤. ��Gn,��i�1�I��3��U��汬W��5zKx�ebv��#u��*:���PaI��_��,\F2���^���<�8p:��K��d�e!n(�n�y�v��M&!�2�?uͻ�㬟rf���|���/�*���?��A��R�g�9\��l7`_���B+��c�hI^�j ���$���|���ԝ�4X���iF�c!=�"����ZɈ�(��s0���@������N�n
��H��G�.�>H�y�������j��a� �������嗡��ݡ�Y�!�oL)�O��� uY�t��/",��L���N�I|j���]#�y���j��אl��o��dRp5�~l�Uo�3l��k��u��G~�i@���Ep�1qy�Fb���+j` D �i�宮M�I��������|���|�2��T��h��QD6U��k���]����U\��J�+��g	�>	hbҡA/RF�N���#1`��\��͓�N#@�1?�>�Э�q���H���p�	iKE}�`���A��z5�ATVAvd��bz�)�����B���2D*���D��+�ى�M�So]#�"9L����b,��z�փ�T_5�5�;O��v�]$>�]u�hz��%�rh��$��d��T�S�ʌJ�z �8J��W[���������Sȹ��A���ZօƁ�����O]"+Ny�Md`aBF���"/�m1�]�>���&�\�Q����c�2'T��QK��5��>c�OIC�N���0�]����jW�E&x�(�\cуO��0����>�N��1sXR�\�:�8D�Yh��0�+�����>��z�	��>�|Z�gȇ�$�㳣\1p�[�:�0��,>[%�v����=M�G}q��Т/&oy|�I^-M��]9,LM
%��g"����$�?1Ș�O�M۹�k	�'p��[wq �7(l#͆�u����JX���˥SGi<J��8��,H�j�?��g���9hړ�D��ʋ����.[��6`(3��V��e:Pe�ї�?hs(Y�©���d'H�|�����<X�Mg,�*�A��y����A���A���Q������MR��'e����N�ѧ�G�[36�XWC�Ve[h�
/��8B�$��p�' c�h.�5�Ul��l?>A���k�3�]X
��B~�/Rj�R1���Zm�I�sˀE�.��G���`�h�ߵ5�����K-\�95k�((�zy��Ѫ����͓��^��4��_}	8G�vI�֖cҋ��l`�<Ϻd�R��B*��5���"jPH��|�ƓBJ��0"opV�1Z��g�yy�����3�ؤ��+�Ɔ��.� ~��ᘮťz���^Q"�]�H]u8��fp��2�p��k����Ε��ɸɹU�d27`�~��"Ǚmc��v%|z�+�J^ݧC�/1�]�HyTף3��=:p�2�r��E��\F��֣3FǗ��2#E���쬉.���q����ߡ��lj�:����ԋ4K���ޤU���H����~;���f�:l��6��A��bO�珣��@���b�p;�����<�c���AC#kX$2g��n��	�-�ه]�>7%�ep$����
�@<��{'���l�:%�H�1bȓ�R����ڧ�/.&��c-� yD�*�A��!�����|������ZĮ nP5�-[[z�/�t���&Gh�������Euwu����n�H>]����h��'*���jGM�Jk�P�)�\Wܮd��M��2�E�0-��+�P2'�ܾ=�E��~W;p$HV��$�o��Z0Kd�E5i��Z]���J��o���=�W{l��7��:�DH,U��7�����c��4j���l�8�1q@p�g|
3���uJ�w��'�%n��j��R�'�Sѧ��,���q���Pj���7x#P�)q�+��W�|\�+���B�Dgl3{���ǣ�GB4�1�X\�sE��^��N�x�v�2l�(�����4�=s��������q2���~�B�jz��8�F(xY6"O�x�_�41yq$���:>7rr��e��6{܊M��2q��Md"
��i縍y��i�PQ�$Y}�(��J��)�,*.�W0r����T�ᶆ�:��n~�&g�g�c�����o���r�қ6��E����T���\��M/W�i�z�D�J�-�|��!�ߍ��/���_��@P
�t2 �u�:ѽ��sN/I�B�+{dGF���9�CIb���KV��NPE^þv�Bt�Պw/H�qE4B�m)T�|���9���7_h@q�e(��nz�OayqL�v�,%�N�3������Bp'=�CF���ǴG	������Xg{?��HG'�5��N�4uԄ]H���u2����hY��'�~Ft/}:�'��k"�P�9�h}�� �?�#[-E�Z�o���c�HN$ʐ��Y]�{F8x$�U5�����!�[�Xl �����Ȳw@�?̥sD��5Wp�S�'����![��@z�z�����BԴ�M�,�P��GуE�0o� 9g�/�(\{L�|�2���zR�|헠Z���d�!oB�H!d��	��	Zw�qa,�?i �Q����ڙ:رċk_-�-Xo��@Gď��ڠ��"�HjFfM��{{�?���./O�&�:�7�G�`Tj�ҀS'!����
~{�7I9|ouV5%�Aڃ�#�a(��)җ����C�"_,�}=��L+���g���wz>gFz�ʦ@x���lc^�S���ݶf����]�D�!\�}gb���
+m�6??$h|��!6n�,O��5��wȍ�jg��z��P[2U�
��㋌U�pr���/$��#N�^0���X�ڢŲ�s�ֳQ}�RWw2���r����a4����vIV��692��f7�m7��"1Q�Ͻ�X��M�a|��Hx�	���]"H�@ 1
X�m�VD���k��v�_�8�{)��̓/n�3���: @������«i��j8C5���p3�O-�~B1�9=��:ZmdFY�{�(`��D��$��B���ⷢI���"EL9�)B�b�#JaPHo�#�A��J���,�`g�v�UYψ���r�n���Y҉.˫9�W¸�=ΐ7��וVz�
�fdOb��B|ܧ��t��<³��ʧV�T�����*�ٰBBH�P���]�j�A�.dv7�"�����~�(����o5qȨ��gbc�C��	AYSp�xp&�*��g���j�(�LG���6�])L�̎��_9��� �Q�IB;�	/��.���&x��d������zzq]�*�8W0#�zqӤ�z-ť�u40����Z�Ko�
�m?t)�U2�8�*"#�ķg4�{��z����LF�P��`^K��������g�!l���`��e(<՘p~�USFK͹N�x��p!;����1lh���ϭ�I����0��� 	�v�>��J�a��՜:��'!������$d[�ro��1����*�L�`_�6G�!O]�������d�!��K�O;&��.�	 �N#iЮқ���ܿ�xp��=�
��:��m�jqP��DHS���Uj��Ȅ��).��xn� ���!���ԧ�@X]�3L0Y�1��R��!�� �"��TP����E��}�~�I�sJu򝐶D 3��¼��}��4Q��Օ��/< H.�O�$)�	J�I�7�2�� ��j.��[7��9����QFm\Q�v�.��R�\"���J��7����V3�������rͪ=j**�is�`q�Ai�t�%c�5�?���gFE�� F�&y*�Q�S��K�m䂎���e���?j��Ơ�A�>�z!ߋ�F-d������L2.<�&_�bM{]��B�T������	7u�b�W�KGz֡�~�4Z'�o������A��3��]�)U��t�C�C��s�x	���)+�4�����ծF�mי�N�E��/��n-wX�Dk���ぅ�B�6T�xIr�e��nZd�X�����k��f/�T���0����P�>{k�3�@1�{(Y�#�$��b�5!�G���FU`[�!(�F\�޺:����q���zE��*OoOp�ȑ	9%��&M���[|}�usD^�$���o�]��>]k���@V����}����a�;c�Ml*��RBֿ�-.�.'�1�oB��ڰ��� �E��N{-��(�b::�O��f���	n����8=�y��8y�lZ�tl�JL+����=�	i�;����tsyE�!�2��G�����x����O���"��6bO�g�L��tn��\�3��!����s�*?�ô}��*s�b�Oc^�	^|�iH��#O�#�����|i�\p%a��z�����y�����UN��F�>+̗�M+\�G��������*Ņ��� pYԐ��G�m?���k1�h��k�5�t�}Ҩ�n�� �����V�)�=@�A�b!'&fmk]��9�N�P6\3����
$���R%Mk�8�H#6�A� 9��V��M�Cc�?��ƀ�/֝.ə�b��RR?XG��Lq5ɿ� ���(�v�z���9'����*\a^�ߗ6�/}h{���p�,�h-�R
C�1m�T�B-�h>�ļ�2ݑJG5)�;�Bꞽz?D�����q���w�^׈�m!
l�o}�Ck`�>�����^�*�OV�InYQ���٘	�g@PIl���$��fMLK$���C�~觖��b��3��E�Y��ب�O��2-w���CH��&
���z�'B)��\�J�a㦣ʉ�k��������9�6q3,�= cl��z��V��/��R�а!���F���?�5B�EA�xM�"@���n�a��eD|$����M0O;�;���CiBɕ��2}Ʊ�L�y���B�1Dȹ�_�գ�̩w�5.�$��p&G/<8�<T�^T�@������$�a�t�' ��J�
�`�|>�1㟝�k�>e���݊]JIc�Bo���\y��*N���er�-����i�b�ډ8�O��&�3�ף��N�t�d�a.T�C�]H�t�s�ks�EV]~;�7s'��7�k�5�WU?��g�@��pӒ�iB�Q>l�e8ʗ����m��
TKLȋ���7h��r�8tX�|N�î��P���ԋ�ӽ�M�ύ5ps�m��-�t*j���&4����FO�ߔ{����~'���6�2��ǼPɜ�����G%~��ܧ(�{�T���
���ë�0뻴�^1�a�|N�%��9T�C�V9=�2�n(#���c��Ek��ҡ�W7�c�b@��
��;t՜�l�A��m-�GtЯ���:��r���,(��3?�3����c}���9D��� ������]����̔���0١5ų�3]�����X]���ݼ_GE�8���V*�J���R�v����آ�x�%�$��*��$O��� �/Q�/@د\��k���jG�i�[ɐ��42�P�s��񯂱��"z|�r3%q���u#Y���幰i���֧�3������h��K��(Ү3��v��"{ ��0,5-.���QH�o�����08���Bt���k4���O�[Y0�d��U[��/6��j^��Ξ? �߫�����Ѯ_{���h$��� G�u��G�m'.>,��Τa��ivD�0���Pu��w��%.5P#��u��FiI渋2�H��=y��4�E�<����L�@ބ���T�J��{EIؼ�2����Zw����rO��L��4������rW-�Y���	feů��{��z��r�0I��␈4�a�vc_���[����n���}�:��<�hd��SI���dd�R�P�b���3ڶ��C��vJ�C{J�W\(M�KwY�t�	��Ǌ�7��\c�j&΂�ƶ��Z(���}���h\=���8T��'#�Tl-]sz�(eշ2�4$��jG�*ֳ�1F����Pޒ�U�W�\�C�T�~��y�r�|#���tֹ��;0���0�ɬO/�iDN�l�� $^@��J���~9��l|u״�r��=oP���	��(��\�����X�Z��w�h�뻃�{�=�J���4o)˾�5�6�kʅ��<��ꬩi;ܔ�)x�/+�r���5�|0}���*Ҁ��4<6ʚ�?��x�cj_��Ub:6�ilR��`�|毙��.4����xk�S��	'p�/�Kzw�~�E���� È�˶fG2;HKx!��s�w�K�/���-�K�w{��
��*[f�]�"�Sd_���s�b_�q�jΚ0�[�C���L�Rn����H��W�6\�Pb s�����^%� emPt\[aD /�b���> �d��
�8g7~R�Z	5��p�������w_6�p*���sfd1��0��bV�ڝI���XfO���w�MQ�L��g�P���&��4%���w�&����@�We��;�]؋���������;۫�ʚA� 8V&��^J��r]Ǔt��Sw�Z+Fƥ~H�ZL��~z(*���	�\�6d���4�����_e���ͺ�g�0k�5�p���.;?�m��;����SL��?I)�J���9?�p%�1�Ut>��3�w�
+���F�P�K&����o�~d�X��Ÿ�5����T@wP�'Ee��J��ዔ}�"�ȔU����w3r)�H:X���Gu����/�{�#��f�mC�o���Z�R��h�����n֩�l�f חҌ�)3��u�TC8�^O�H^�������i&_и#�%+�s�s;��sh��R3l�'��'��άl����\���a�~/H�ZPU����f��)sr�Yk��f,_�/�~i��Z�6o��w�uR,強]-û�c�P���1�("���ֺ�/h�Z$����l@��5Wya���}B�"�au0�%Za��;� �P�J�;�K[2�[�]��\^4�zE�Nf8R|Ƙ[KH<����ORe�ݎ;sk���BM�@�X�> �5�A@��e�|h�Hؒ%�)���y�i��p�Bz2Z� 0�\��z)���i���W+�Ƈ�EBf`fo��mm���;E�	D���U���þ��k	�=����k�Q�1���u2�\gw&��VI�E�m��u_ȳ���n�`�~"���>��?�i�E��Yp߳���&u���?n�
`F{u���dI�ֽb�m�i�ْm����糒��oV쯌�(��b8PF�X���^R��R�^Ymǒ��؍�ߜL0g���~V�;�/��@=/-��s��t�N��"�x7�#D�^g��\E6��l$��j��4��ޛ �/𧅽��j��{�a�׷*2l/�)r0P��~-�<�]8C���9W�#��$����*��eM�.$�W��o۬VF����Ѝ���3���H��#&>�����s,�\�H�ݺ�2���2�T��6�*Zz:N�Ԓ;��K�fƠ��Qxվ��x&V���~�'���E�/Ƃ^4�z�S{T�piFk���M��b2/���K֔ ��I`��S�kN�C}�ZL����o˕Mi��k�Š��:eN�'}�L��GO7m`�BxH��C
*@P}��NTa����+tt3��(�˭F�ҽ����;�۬Y�N��@l*���ɭ�L���K��5�ϴ�o�؝ˎ�`��t�֠���ǉ2�	�7��7�������QBm�n�J[����K�xh*�2�� �U��P� ə6s�����^"+`��i)H
�p���w���O�)��H�l����`�j&�M/��AX��vi�V�)t�p������6���]F��䁲 T�]p6*��T�L\��5��V߳����)��=����?��(�bIL�%��X�Ho��J��%>[�ٶ̒�ՙ7���#~�>��3�s�[�#5�9"���E'������x���m{��8����<������t�P���L6��Y�n����j(�թ�
�I[�X,�JG35�ׂ�I�V}�̡2�����-1�~������������tʮV�^3�\�	�T������6�o����h�5�\��0ޏ,��$�+cѵt��	��B������O���O�<C:�0�}
�G����ǻ-��º���-��oB/��F�o���������M�nS(IHd����C�Y~[��η�T�`gܬBF=ۭ_��,d��0Q�V���22�̗��P�'(�8:��Kx���oӿ4��P$@��ݡ��v���\�8���c���j+�U2���eD'e����0�R�/�?m�" �rv2�JN4�J�B_8s|;��߷זYF���و��9�)��#���b��d��Ruw�w��ے��V��_y%g�����JO_��O̵���	!v��CM�-��3RgL?����U9N�����BB��*��>�i&��\e�~":��J����U�D�&����+(S�׫� �f�Eդ��o���!��� [��I$TT;�n�L��aJ,zz���vm��Ϩ�2A��`�;u4�3�Ԉ����j�&Z��3�'�y�e�Q�i�g�����`��&�k�@SS���w�,bxTγ~&���u��Ki} �v��F��T+U:�?C"����)WAA�|��N�}~�֤��	�MkCf5&��mB�M�Δ��@A���p�:Fn�j��f6`׸��լ}lt����L �z�73���b����B����7��������YYY��r��p��N�c"q�hG�da��_l�m�d�Z��sK��>NL.��6�]��=���H���2̖����|� ��Bx��i�1�Vx�-�=AOƳ︇�l��`>�S��?�h2<d��)�9E:"ʪY��]zW�
[1����d�̎	k<f�#-���4�����|�I<x���BA<��A�K(Xt�v^╹ V��)�,��λ�Zt�J�j�9)��S-���Z�YXݗ��IVϲDE�K�wT/����!��HF�w@}�ּH�P���4�%v���%i� �95%�������?�*X�h��M�C����[)����D�f���^��̰t��BJ��A�$��}��rM�!P�^����l��M��=���1���F�͓B����}K�ml�����]���
������. o���āf��?'�F˘|�q�>8�[���u
�A�H�	��$tQ�o��*�9��a��Tљ8%��#O����'�gzK;����K.�`�sz{�d��EH ��I>^�y*�����	�o����6�t[��s�T�a�_9���@��+(?�2�,��V!�%�X���:��n�q�^ɼ(Ym�� ���Ҋ�wy�2��{x�;8����߹��Q�ؽp�[��J��2eAP�ωg�S�M�=��ٟz�lbPz �
�����P3(.�E�l�S�,�̣�[L.���x�cԼm0fD���~{e�B�)����Y���ё����XJ��*�KM��(��tsci4:(3T�^n4����K�NrA;wz�Rck&p�J���e�˶/��9���E�U�mx�8R��E�z��l���48޾�e`�%�|�����$��N[L����?��S�?j��/�$�LL��5O��U�1�o�Ou�&�Een4��f�g���x��@a�q����\l��ؓ��:��@v1���gB�q���E4ӝ����&�~�=���
ȅ,m����)ĠUT�v�R�M���?�eլ���ô��l�ƓH
f�D5u��<�k��|����VZ% Nm�9dC�H#��� ��/�������������=�ޗ-��G�����ޭ]Z�vع|�/�5�	�w����2cݬ��O���S:�h�N"s�ٗ�}}�EJ��,h�Q�Ln�b1V�����(r-���4���Cʞ��t8$�c~��8J������a���8�P�4�%0a[w��[����>ի�vPf��Ӗp���p���Ւ���&�#��(��1 E-l�G�z��R��V-?la�KR�T��Eȫ-���&�j]cY�h��'K���8�_m��.S�n�#�B�/>�IW%�Nt�s�]g9�b(�Ś/E@�@U�^�M�FN"ب)t5���Y.��e�֯�������]I�Ia���mt��±��tlM/���-��c(��lfB�����w �����8O�Yx�L"���� `f�T\>�M&���Z�ng��#���&�]^7`�,|�E��0e�;����>�# �֢K��韺�w1��|^S��8-V��͒�{���%�����Č=���˛A�
h3G�����q����Q�*'m��!�����I�\%���Qs�!j�lr���s�� ,�C��[B�BH/���ü���"՞�i�>(_���B<^]t	��5lI�k���Q[K8���],%�)��0�d�`q�mK�HL����p�q��(�_�o��;�R�1�h�McU6�~S���;��We��+G:9��� ��6�"D�%c;���Se�;�A1V9{�q�  �:	ĩc��t�_�5s˅���:���/�F�IH��.C^�V�Ѵ���{������,���r�e02�t-#�����Z{�ޔ���g�¾�{���f
R��; ���J�}Qv^hLcr�1��6����$��1 ��K>=1�mef�_���ԣ�t��j�]���{�p�Xx�p;�l�>���6?8<6bZ}���> ��a=B�eʩ�h��ŕj��&#��Hx��=�qn|��U���=���ו�OaJD�y0�`��J�����#�/��2��E.qn���^�_��>�D�-��\��#�����Y��tV����9�-�IT(_kN��R���e�T_�J�uw߭��&Brܥ)c%!���F�q����;߼����Yr��~N�?c)-
�#(�(	p��L���˻]c%Ν�z�seS���'}[f:�̉�|��Ӵ0�C8��!*�Os%�4w;�wƟc�3L&�{���k_@Y��r&��k|$���:U�=��hT����ڲ-��6
�_��ݸa��F���u��H쯘�0��?��/��a�u���
�Ϲ�,�ӳ`��La��W�m�ݡ	�a���%Nb�+0���`wɗ��v���)���1FsȽ��"L�F��g
��f��+�abEj����.�LC"!���r���w��h�=�������!�����-�m��>e$��ڻ��i�)��!c��7�(��n֡��=
�#��vp c��e��N#"O�wA�5׸�:�1;G�ZY��o�vf,ĚW��-oV���d"J����Q蠩�/�qQd�ȵo���E��o���j�����t	�:�8�՚�R�b�o��t9�c
Z�Vo���\��p��*�~��b,V�z���� ,�7���EL����z�^�&�R������;hږ��qs,��8I���ךΙ���B�WXmV�㥹�0N*`������΃����͑ߤw)�~"R���C8��G`��С%��C�P�����\it.���/�����O%λ��@x��vƖ�H�5Μ���
e�P<��q���?���]N�l���D��:~ٴ����Ζl����A�r��`Y�W)QX�"��lr�E5ғ��/��5�R��R�vo�&�F��Xh-���gٍ���/���BG�3��q4���ۄ�+�z�l��pЗ0��J,Կ��������Tv��Tw=I����˷[ac	M�ܡ*'��Ƀ P��u~<v7�-۪O� ~�c�'��W��L`�k5��RY���k%�pua<=���Ox ]|�{}a�%]@o�Жn�%��E��ϩN���\^[%����z���P|���E9�
�P�Ҝ����Y`R7�YDN�?]oG@���R7<��f�g/���Z� 4��1��g��4���=0Ҏ���g_�>�E�=�s��Ti��\nr9̀[��2�x�A���{؊�O�\�?���F,��ѽ�ih�RГ����0��y�{���.F��^-��S'5��P���G�T�����
H%qNeQ��Ch�[�J4|��3;��0}�0j��x�襝/a3�gm�AW�g��,|�sG����d���JL�+��&�.l��L��� ��J&�¤�o��"ja�I�;j���eqm���j�oS��+P���I�I��=�O���L�OT�X7K�Uv��DobD��>8�;X��,9��f��/�4�Rg!�t�+�I���pPX�����y����������{� 7�ni�y��w��h����pQ���pZ�(���§�$�lK,yƧ�hl��<�X�V���sk���v���c=���q�c1�R�4
���(.a��!%��Ϊ��"�;>r=���hg�0���������獂�#�나Y$�Y6��L��{��2�^�2��x
�ر�>�j>n\u^�'%���]­ǒ���m8�p㾹��T���OP�3�(�^\oT��������0�,��u�/�i�K��W�%ZR�zƮ�\��Ku�ellwDPQ����8���ѡ��T�w�۰�[���ܼ���w�ت�V��vT�Y���3�6�ް��x\��klS״�h��K�{�EF`Mqh����6����	Ҵ�hV��"�t^f�V�1Y��ѳ���dH��CZ���o� D��C�6�DOs���~����0$}���ئ@��{`�x��@Ŧ��xn.�v|��&�^ƣ�d���bYQ�I%ີ��=Lt+X��^��ҋ��X?�Akz�����6��s���%��47�ɚ�Ɏ�L9� &�3/1��	���|f���6P���yv�Qb=�X�L��it��#l{2�'���y]��g5,7[>�-w��vm�z $�A�E�Q&A&>�80 �2�-x�u�����$��21�k��x���Ȥ���T�o	�Z� ��u��K[��cHR��<9����})�N��dt[���T��*&��K\��0�_u�,y�A��\P�g*�Wm���	��3g4��V�sYB�>�\�{j_V�I���+�Žو��A(E��%R+�|�~�QT��8�ґ�@+A�MMq�"��׳R[r��n�Nj�3}Ǟ�c?JM����c������p����
�H,�ܼ�k��5nE�e�)?�5����o����[�P.�d��(
vH�n��<��\�gFE^��B��/�+#�@p��9��$�c) D�}�Ӷ?ҭ��ή=��#[yÎ{{��)�9lu�+����Wzٲ��������k5�	�����(�+����A��27�܈������L�М�@�-���m5� Ĺ5q\�Mdjo��FA/�xs�V��4Ӯ�ga}�2�X���'r�r@#3ݫxW>H^����gGCM��B�_m�h��D�������~��8�RWD:���i8�攒O1w�����o.Ja`�ۗ~	������yU�!�J��ýN�!��GoÅ	`d��/���25-�>��"�2&(nP2�h�m������M���9쫺O�������t�v���?]�۹���L��!"W��˜SH\��%�q�1���uީG��$���+K��G�����:G1��hib�TGq��^��߰,09���(4�$�@����}�o�XK����⹯H�VT;�z���	nwF�JU��7��ȿ
��K-X�:f���[y:���?<�g��o9�x�7��R��".��m��V?�����Ki�|OQ�-P8���U�`T'��`+W4�hfrT���z�b��ln�H�/��.��`P�[L��W>�����r���o�~p�e�?c��*����&>R��]��8O�S��ԯؑ��`���;�@iO
�[��C��q�oilG�� 9$*�u5h�a�=��|v��C؇*0�T�Z��{C���*�Ӯha��s���s�c��c�Ԡd4׷�ww@�{歹X���}Z줐�'��`���ils�B����J&�� ���k��ښf^��*n����oZ;��M��~����`z�����×��pB}R�V��8+~S���Dz�m�hx�ʙ��bBU�8#ͼ�ҳL E�6;/� }jGU)#�b���٘#�n��X������L��	�����A��MH/Kp����}Ԥ����TG�w	*5��t�#�~1�,y�뫹γ��6��m�m��j>B���W�ǌ!ze*���<���ލs<����I�S��7{����S�l����SS�έ�[+e(��'�&�Ģ��Խ������%�MMCN����4��ڋ�9�ot��(z,�;m��Avv����D���;���[��ǑV�VVMSS����b�~zT!��$�=$��l�=m��A<�Lf!�
D�s��Wy4���	D[��������v|u�L5[��p �|Q�fr��h�XI!��sM���P8�D7+禲���a�g���LqR�T�q�� �6��9sG��C�d����<�:Dƻ�MZi3�T�\sc����"��Vb��n��F�iκ44��Gfi���MN����8:M��U�mP�(TX|_/��`0�'%'Y����)�&���~�
r4��BB"�γ�+VT8�̮ӛ�*}��B��GL��d��Q�}Wu��i*�MNc/�$$H�������1���9��Á�6�+�C��u�=�����ȶW"g�\�H�ZדR�)E�젷(��>*5���Ş��M<�.�uqF�n�)��hq��"I�,6�����1�ksӥۛ5��;�,^�9G�l��*!@�\[�{����T�XUx`�7�:WN�zHT��/u�P����
H&rY��r����N3�դ(���l�O��#4��hh��IV�*��'��[-�Fz�QZjxR���E���DҎ�oP��$aS��L�#Sޞ 3g���m�+&���:QH�KS���������~)#^<:�_�,��..5�#�J`!�	Z/rP�����/ R���1��x�rպ�V�~=��:"N7&V���O���Un���×S�1�:ͪѨTFE�=�C��X��p�a!�]e`��r����ꈰqQ$c�[�V�j�zEJ�q<��M��hG!�������u�2���g�:�C��inI��Pak�c[Ñ"�ǯV��"��"$L�GnM��EʖՎ��"��w�P3� �)~uz�8�_���&�����x�~\��$�"О+�KTy���8.gOB��&್S�`&3P��:�#=�0\V��>�B~ѯ����k��2��c�l2�ޢIA�]��W�����o���ڨ��������h�!���?(�wn����9_Jբ+yf�0o�!�A	�4F��]�R��t����֎���!�*������~ˬt||����ܸꊕ Z�l�DP%���u�� �"Z(A��E�ƈʚQu1���G��|�d��\����ӭ�	��y�7s�d%쬑��R��O���T\y$%�%@��z j�D�ǣ��k��V�1�@�+n��筷��9=��~�w|؏���ǅ)\x:�]/�2�_9�x�JA_�]��E�D5q��v�i�)�G�[W/���{��Ѩ�Ky�q�³�Ѭ5��c��qJ�X^�Cdl6b����m�߬�~���=EH?����&��qi�:�X\�ka���o��J��~�"oo7'�> OX�~���� �2*`�I5���>a�}�$ b���<m�b�hmT��ʿ��[iN���'*J����;�]jӺ̛L���/g<$�{p��U��۸�i�3��+f��L�YE���vuI����^ځ'�+�X�ѢiZ���zg��\��������"Ł�{�X��օ&�	^����cͣ�%��:Ip-C�J�o�������n��2!̃ų�|*&NXaz��/%�j���S��i>���aN� �!.�2a�a�l�K�p������4��,"͡��7�p�s�#W�D�_Y�j!XOx�7E9�On�� `�Ѐ��m��bXXc����夯����-E����wq��ܢ9��ڊ�e�{����j��NwE���e�q'�M��Ց�!���$�[�Ě?,���N�@�3���'v�nV`�/0&�����5Α>y]K���{�Be@�*�Zf��{H]J�]��?O�~5�w�ڎ�:���G,="���eKM%�Uڦ3�jU!|"��O��+?��u�tS��{=��+z��ŉ��xj/���������6�p��B%�w[ũ�-�&8�2��#7>�򰄘r�x|��'0 �r�r�%�U7ٵ񩆗[�%��f�&
a����3&0��v2p��˖<�. {X�~��Ɍp��4���T���^?,�znu���ԇ̢�;�$�,��3+���=pc�s�T�z�ppq�I�5+Q��˷� ^��f�x�*���.��wE:{������%I�����G��
�@T0l���� �a|�]F��q}��1���)>l`��٧��"!:=,9����t=�q����#��Y�r� l%u�[��o���3�ܷ�+�r"A�5��J�����[��>�b0}#��Ig&+R���x�;wJ��4��%/�l%'����ӰJ��Yt;(�?Ǆ�i.�RĀl�R0�X�Ҥ�)�Pnٍ"�!��qx"eVZ�8~wH=7$�^�9��Xx6]��R�g'�����m��%X�_3�o�ɪ���k����,=��h�G�LII�&)�Xb����.������h�8{v�
�w��թ#C��b���H�E��~��F��J����[�4�YG���s G�E��Yфi��[��"�M�G7$X�r�k/�_�'b��s$��W�,%�6
��n������vu^�)~�uP�"e�þ٦��x��g�+X	!��Y�6�َ�s=���-vD>H�0M�� ���t ��f�Z|8ݥ�Cc.��к bk�^�d�WtQ�1���K������,����6��+^y���eg7T���oM��۹��FJ]8�d;���m�2�u�Eg��>�[@4�ఴ�2p�`�x��5��13"�x�*�'Y���[ŉ�K���|T�%�����
�Z� �ڨ����SZ~�Ǉ�����̦�~b>A���P�U *Q���ן����?�j��d:�pJ�P�/vY}��,�P�y���r ~�ji��46z>����k��0�b�x+��H2^�4��_̥�Y�[�mm=��5Ō�h����Q��^D�B������a��e�����{y�c�Kϼ������q����-ao,=(��z��k�1x-�,����E��^�r Yt�1�*#	�#-G�3?�D��x�>�e��@���1M���V?x&���c`p�q�,�qK:����A�~fY�2���ʜ2]7I�`@�ZD�N+��!c�	���2p��D&g�N�K�A<�F4:����j5ט3�·�u�ж ��e)�X
��_�s����v� �ͅ �W�":k�g���f�r����Ve�����%�)}$���_,#/��*�n���R��6#y{����>�7��o��*Ue_`QK*aQ����cW���C�K}sA
��Z�
Z2�dEmF�՟R�bh��A��-��+d�B��I�Y�A����9�v��J�vG��H��]�Gi9!w
�$	��K������+c _e�;���%!�D�]H�4Spo�bA>��Qxf�h��y�W�>����������0L�MG�UOQ�>B�*�c����@�������3��O�a�h,�M�m��(6��̤[���:�1mqf�ZO�;��p1�%v��V�ʐ�.W	��{�l�4����y�>�s�G'9fo4�*�M@\0��o�}���>�D21�[ȑ�y����'x��s�|���M�ތ˥a�0J"�c��l��cG�F��st��x)iyZ�uk?�����7w(\�V�+��~L��匉�l���.	��9����EⲔp���q9��g������3���T���"
��5j5�M�Te�B6��Ea�@���W�=�&}Y�q���ԯpF��X�eQ���x�?�Y&�9���i�r�iǛ�����E� �d��N�a��O��ɉ=g�M���~�&<=t�j�+y\��c��������P@H��˩�WK׮������wU�0���B&����j&�4�ʐ�_�1J@��lS>)��cDe7�p��s�#�<4!فgF��2�Xvv;_P�����ݖ] �1U�um�aX�0�`�v����/z�����c
��R����D��S_��_�~jX;�COhF����cX�U9O��!��O��[=/�#�
h�ه���`6BF=`�T����o�A���Wgw�7�
� S��(�LʼQBn^|Ƴ	��k���sG�@oU��Ãѧm��;0���U���.%�D �鵮B2W�u>���R9q�?�Y��Fߒ��v�p4�&9�~�!� .�4*8�e):����ˤ58��?�-A��^޽-`V "�V�M7���\׶�m�3d1c�'�+�@A�H������0\�y�)��'TSW�R˙���9)z�8�ɨE�5������)'��/�Y�j�;ؼ�J����i�`쿯L/-;~Ƚ�x�4m�5C��r5�jܭa:v�c(J�(�:7(�3'����q�7Z�`�c9Rn�P��������'H�5�hV�Ce?�.�"L���~�� ܍��mw�6�p�v&����Y�Xϐ`R��بh�0�n#�ຫ[º0��O��t��BwK����U�c��IئpK��#�I<3�]ݼ�-�-��j������E�
�:���L�}�4�W,�L��g�3�u7�'�n�zZO��HW�m�Y<���8n��#��r���n�J�B���jV�A��L���p�D�4��3�t��S"�>���#nQ�-XDe� Op�e����\M�S5�ǰgqS�6�.���v�j���7v�F�B�k�ǈ=�&$�+���G�8s������sy���d?����:��v���l�~�yd�+���乕C��:��D8%��֙q�m���-���KB�ϬF�A�D����Sށ��1CĪ>��#>�`N�`tz�Wj�e�0�D7ǰoK����=I�p�0K�R%(rJ��kiOے���(����>�;�����īB �*����j����XlxVHYEB    a24d    4340��.^[<����e��z{���r�(����tgfB���/�m�<��׮�>�xգ)t��p"G���W.و�f�u��M}-�Y%�H`� �6�@9!`��-�Hz�<܎�����p��u���7E�C{Y�
k��Qk�|!@���u����b簐��BA R�����x�,3$�yDɣ�0 ���	1[�e�ϻԐNd�-��sa��R�c�7V�	\��z|�B�LM�����X<C̙m.E�-=H�e�41�_X5�_r�3����G(&���MU�ʄ��m��dxY(���TLAy���,D�
�p�/�-؅�~Ԑ7<��_��}�����.,�� #��}���f��`�=X��(#�z��hظ��zKMo��*�����\��Iv
����o�6��V����W���J�ڜ��OT� iH�3k/0��1oP������'\{�7�<_*������[׉��߭?�B�h�2��F�=�����K��z������'��F5��/�xg;���:����.�f��T��A8\8Mp@�ˉ�jV��@�C�6���>�wન�TG�T^䛃�3}.�EI1W��iu�/_#L�����w5nY�>��4����3H�ʇ4&������Ǉ���5�����}��g� �>���%t37$k�wO� K\$<�2�W��NF57�åa��pUB}L�3�.]	 >S� ���:��v֮���ub��wl9�ba:�e�W����~���P�oV?@մ�-Ϲ��:&AJ�E,��8��?�0��r+^ �C/�u� qNꃈ�|`s%`ɲ_�� ���V��,�j4U^��?x~]����g�zg��V�^���4����F<i�=��Փu�+TJ1�=^V�.�谍MY�G���"ɽ|7�u��w��+-ڬ���-(Ӓ���Tl���>���W���4�46��:ʞf�#�PΩ��p(9QX��8c$�>�yI(��/z!������S_�Y��R���.z�ā��O��{���Z���Z�U3�=�80f[��}�0]/��l�sS!�\٥%aOm�ζZ:�ūZ,��"��x	A���P
V�l���[��T���82��$6�Mj�����J��1��hi#3��CW�gS�n_*zL1���yF	]ƣ! ��&�"�	y�`��KY�`�����!L,e@�����08γ�߆��{V��5��Z��o��D �*�L�O�r��o��'2�;�Y�|�{������ْ���ji�;GPG���T��T����d��V�}a�����ۡq,ԡPԐOG�X��f�{��:YQ��2�7*�N<>C*�*�jwx5Jf���L���OF���,�}�Bu'���V�wҿ�U�ZA�k���W疇���ٙd�dk.e�}件���gΒ'�jv�5r/(� �-��Ĳ�-��xdY��,Tt����0�R����w��s+�5��h�$��G�G}t4��]�0�R����H2�������6玉���\�x;{�$z@��4P�3�d�Ri����j�0�.��:Y�&��i�
&�X(����~��na'|��>�[�Eu��T��F¢C��{�>�_�t�\⢐t�D�x��X��?s�),浪���[�{K��CS�t9ߑ_s������.^�v~˜�.���n�<H:��%���0��#<�{z��0�xl�0�5!��F�,�{m?jt�	�cNf��Jb!"� �`Z`�ewa�}��<�'�9���(UYp�����M��tA�
���|�d��ㆪ���#�K+]�RO�B{��>/j��_��l���.��h����gI�1/��WO�1�:�_�SQ*�s�,��� 4D��4]l��H�J:��9@;`��{�蚚�o�X>5���2�D� �=XVt������љTV�$Q��+U�-��͏���.l9�ٴg���c|�@ym�hJ�hZ�H3�=��"1>�3���\��2\j�M��W]���y*�^(�N��P��w1���2�d��ה��[����-V$V��?c.J(C��IK����F���{�*�����T_^�{f]9l�p^���Y�Lk�NuucD�.
��ޞ��?���}T>�ՂI�?`�e%L׊�ƄMcf��cv9\�-i@Do����Sz�<؋�{L�=!�zB��m��sn�]��Q/S�p0;�7V{G#	T��Uw�>��./����a��4��oV�X�^2�W�	_]�@����]��_��bX_����NS�pvh�n
���÷�����1-�q6ե����L0�#�ǃ�]%����E'���D)��t6��hhQ���� �*6|�����?[��&�30����SHm&�˻-2/�(���r{�D8p(x�]l�j�𦧔ސxx�
=y#L�u��~�@cN ���K�>�LU�[�[��f����th�5?�<�x"���D:N�k����2ϻ�H�v�K_��:MT;�4���Ȕ���5���7ĸ;X8�a����-��ơ� �����$CY�a�=mo�I~Xg�.cіv�����]�P��yx`��lm�����`����
vg�i�z���u��8��(м�S4a��I�]/����]*R��9Y��n��F�<@��̼�Zֲg�(2� M��dds���*���t���@N$^�(��џ�p�n4gCe���h%��l)��%~]����j��4������m�P�q�6�4����U�`X�Fmte��P�F�U�޷��T[Nܒ���Y��<y�œ�;&G۬ �*o�
-K#�k�����hs��*�����0��sK�S���Q3�b	[Z�rE����Lq"�rb�:�F]�]dm��WG�V�I�B��%�C� �QWw&�^/�ͧ������7q������%�6�������"ڌ��B���ʎ��[U�g&\*\�6A���:#�XA�⮸��j+��i>hZ����1��6%�r��j{����</J;
�L�1�L�� �����DVGE4ԂơU�5I�0"[;��Չ�7�!0�Xۂ"E��}��J�+8���o.Ŷ��H>q�X�a��3�����ǀHy��n���
��ɜ�J���<�+<���ˏ�Vrb�t��
(d�[�5��%��N�Mн�Ѯ9�9^
ֆ-�E�qm�s[M澐R��y�L#�\������������#�I_ %Q8�������;ߺ��^����hχ�ɭ֥�<�7�8�,�lSd̮���}����k ����V�>�[xo�����Ky�՚zR����F�߁�T}7�e
�4F�5�tE�'q䡾�j �ڜ����z���;��ٺ&t~� ב���'�[���P��ުL�g7�t0*�Q���}]�F��$��^�7���U�#�7;�`�����a�i?��]ϰ�t�����Z�n�},��!Z�g>��r�ȴ��so^� &W��	@N)i��E�$4��j!r.yR��9ho���2 ��J(��9�\-n�WW͉���F�Ac�I�y�J挪c�b]��q�ny�����r����o��A�;��ˮ����W�m�p���BֳT~��y�����tL��ձ��)��)�vbwX�*J|�7��/��i"��O,�|�K?:L����EtP�4e�}�9�*�K�f��;NŜ�)�Ң�oW���Z���(�-`�?��F.�h
�uYp�^w���<�$e�텾"8I���/'�/�Mӝ-n7.��!kI�-I ��'��=��ݤ.a�5-õ�{�#�%�עVYd�M�LrQWߤ�}��@A�O)sQd�:�l����t٣1�:��O�d�Y^��Hy��{f �5�m[4Q@��-JU~�U����P3�, ����C8��r��V=t��ackKl �7��hl�Y��:��Y�Q �澒޶���^��7҉���>�2�t0~������B�ẹ�	X��g7[ȭ���P�Nv�I��7]��
�M�n��4�I	'+3��ۣ�N<�]�t�`�[�� ��8�Hy�$�\�%k.��ݒ0�c`�5�D���DQpj�h�K�}d�P�mC3fa�%��]�5}'�*�m���q̛�h���U�����1�<�Ti@�� 3!#]��L'lN���w8_UF1��5/ ���0�����>�MEOU�� uWr���U��!%�D�k-tY=2̑Pm��A�Z�q��y�T�R!_�)��}�A���9���.
�gā�OHz�O��|�=N��?߄W:��U�Z�3/��o����Q��7�͊J�|�><���j	҄�:(�bgK6&u�`b���\���j�hr�{Z�B��ÿ*���"�5�vn���m	7�	lm���O�a��J�q�h�h �=�2� ���q�Kݝ��m��E�g��a�-J�Ԭ�`��,�W������B��a%BE�L�7� ��Z�eq/����
�A�8������'5Ѝy�Xr�~�|bg��j�!_
i�y.���g���$�Z�����鋤9��׷�nS_��2��O�R%��������SA�<��*�AM���*i�'�"6q	۩��h�'���hP�����P�U���)��v��q���[��\�,����d�ve4	P��^�u�<�G�����"S����V�'P�T���nw�Kk�v���kE^�%	���rh�@�B���(~�+}0�f'�6&��i����/!�1e������fA����&�nM|�h�䁻�{Kܿ��8��b�(�K'p_���Cl�݈EEtGw?I�����<�x�f�&�¡qU��೺�U���x0��o:1csfog�,@Ө�'���t�g�)?�#v=jd)��0���H	�?�SK�y+[�Qt?Y묘�u��E�D �ª����յ�Ъ|�0���ڐ���/�nK��ѐiQ�z��3,�k+Yժ�:j���v�oљ �+��	��>��K�:#��¡J�A)7˗9+ 1nM������
-v�pr���X��LQm�8��4�ɛZ�h#��tN�����"	m���Lܥ�]ү^v��ݣ����M"��>,��g�#�8�T��K\MT���V؇&�N��|�V���!��|�"k�=g�_�U���nb�V6���ŎAN�H;䇲�AB��/t��J;�dえ���t�ԠX����ΰǜn�˅�rm��1f���T⧹�����POE�RyR�j]o�2�0�X��G1X�c��
�c�!MU�(k�K\�>s�|��ҍ�'�}�Vy��W�kn��+	#
�h��H���Wh���S���1����yy �=��&���K�����{Ux" ��sflYb���>2�����Q�]0.���:�J���\Pb9�u���X����3�Wͩ՜�MD�q�H�h��=��v�)��ļ����l��,/�_�*�i�Du�i�$�\�%����P���i�z���<��\����0�VzX�\���q�b��6sוȟ>�A\���Ƞw+a`�۝�	��1[u�_"����q����g�{��f^��kf~��f��tNx�V(�>!�.�3��Q2�D�&�I�]	��0L�B�,3��+s�F�v���I	9m�$��:�b��%"�F�?�b)�fhXcy�����H��:�+g; �t�Y3��J���q��+�pؽ<�#���mW�|�s�3ݱ��G�9�D��R�,ϜlT���K�B���l��]-P�7f�u��yK׌u;�H[�G2Ñf�;��L��ы����H$��)�<}��:;,_}c���A��W4����U"J!��%��?V��H�4�r�'��3ȍ�Ъ=���r� ��*t���μj����?SjLpB[�P��.��e��1���s.��7�L�Ek[��c��r�b��L]��Bn]�>�%D�$f�Kؖn�3���q{�xcJ9C��'�m�U��N��r �@>�';9*��Sv1U9��p:q&�Qp�'�=��� ��_R&,a�'2ᝎڳ�(
0����\�&���&�e���}��	�X�~�=Z^�b6Kz���T�K���m�z{L�����܅]a�|M�,�5V���s��&s�r��X�$�Kv����?��#T1�פk>,;��5q�nS��.�>24�P&3��͆N��۷��M�mq�` �)���3D��Ǣ0B��?�eQ�4��Z� 
=3�`y�R����d�M������_Q��M��0R�(w,��Y���b��E��F_v(1go=��H$�o�lF�(�'�P�1*�w|o��U���i+�U�����P5�}�����z�T�$����r�S?��� ��.I�8#�h@%�_���a���U��E.C����
��0󀉢F���[�6�Pރy^�5���rxȷ`�/1���ɝ�'��Xq�tJ�i3E[�]W��W��3.�k��C�;A�i��A��a���oPaF�
��?�^���F�0�ݚ��$�܎�5o�'��[r����y����+���~�}w��'g����
�vO�'U��Г�A@ri���!�c�fx���O�\q'[�$�7�ހ���T��d�W^�q��,�w%>mG?�F�YS��A��L�[�PHK�^��ԇeS�]�#^ǓX���k����;+�;����:K����
�R�X�䎧��#j���W�Z�1bŲ��#W��$�<ȫp���*��D��.T!�f��2wUn��s3�����ۗP��B�#jяV���#��H�@��Qɚ�S��ϰIN����)!�ߒ�MM���iT�=��*��QY�k���nVJA�I<Ka85�����~�*�A底�Om?�� �0�v��/!T��b��M�Y��f��`�uXYm]�6�JG�w�*m��l�ȍ[U�+�z��`��ز�	���3���F5u�@�^/,V�V5{.˴�ز%���G@4��f;�������j{u�l_>�rAD"0g=+��_(Ht��w�h��^ͯ���Ox[�,���8��:M��۩ ^�$��C)�7l�,���x[�G�$�2q.d��dMx�0?<��4��r ���qv{�W,v2��o��#W��)�]K�{� ���'�m����\�\�.<�+��C��M��7d:&������GЁ�7�m�ύ�F����� [k}{��@K3�ٓ\'9雬oW�i�{a�e���p�JM�����kW>#�ۉȚm�?��/��#֘�]��XN������Zi(a��
�;b�o9�d	ł�Zl@ym��4��Zm�O]�7����ԯ, ^#Of�o,�7�$��Ic��4xƤ�,���`�ip��"Oƻ$ ��$!ʈf}ÝD�x�%s�p0a�K�;~(��fn�:N�� �W�5�6W��	U?te��E�Qw��	��7G��Χ�8y�N��%޳�V��e� �ٜÆ��e<,��SY������M�<�bP���W��}KS�,1Y��]e~4|����>�sg����V��ɞ�U�3vO�А�vX40� c��]fOR����0�1<��cW���@�P*qq�g_`��^ܺ�frU�k'r�����$zo��Cdf����-�8�+,�,�UA(�A,u��of-+�a;X��)�^茐�ɝ�7t����õ�-f�*�Y��r�G�Y��D�#�O	��̀��Ѐ$�u��t�ݡd=�-aG��[m�2$����^��\A��؛E��X)q�8}�n��h�o�.�'�� �I\F^��!&@ ��3�@u����M�<���5D�քb�^����/Yo�R��٭NA�~���W,�}� pV��E_N�}�@�.h(p�r5B딩x��M�X�t�+�<C�F�cD�B\��ft3.?{n8���G=^��.�vI���I ����h�!`<�&"�ă��=1b�6:�4���`�N��=pMkKǌ�a<@u�/%��(kC��s���"G[���k .��|��n<��wm�b��m�W�M���[6ݖ�Nyaq֠���J+���2 }���D�<�ѫ�!FZs�67d�n����/*���kD8%�A���-,%�b��Z���P�Ϳ�er�|_��k~����1,��@���Ee����Hj����Պ��T�}Xp�����Jw�ɂO�|�Ѓd���r����T:K�W�.�6����(��Y��-v0��-9�iO�O��I�T����)8� �z��L�R*_��W�� �QX0?�d������8�,џ�9�B�����
�3�)����=E�d^;�d�� �ޘ�E��O�h"��ڷ
�7�5�q���GD�z�{�L�H�1�X��轂�H+eL~�r��)��!IS:W; ����������O��u�`���p��'L�i�������8���*��q�O��2n�1O�Ym� �)m��
-�̚B�i�T���ԛ��ݣ+��L؂@k�l#�p~���E��~ ��}��\q\� D�@�.��c7'<v���=
���5k����$���|�{WyW�/i�B��kj҈;O<7epZ'2-�%t*e�2(�V{����`�-� !xj���C�Qa/�p��C����m�Y���D����-�d�a N�&��ӱ������(u�O��$����3�}�������#d� �}������6A,���u����ŗ��qx����A���� �� D���Ws��ˌO�r�ET��[$�,�b�p_fh]����T��y0Q��D��?���d��c��Ŭ�����W\CBT��1�J,��־���p������Vժ�D����'9��,5	C���IT��L 9�t���NT��-�=�N�6O2�c�2~Z�W��6��b��W�Ԃ�� ��_��Fs����C��o�R ��,\���	�l�,�w�X-h�c�I�Im�k��_�<�{��W%KZ������[XZ�]^$��4�bT'���S�74�]ʘ�a�̉k۳M�*~�Y}�̈́�o�o�Z������m��%�9�>T�?g�oJ��C:��O��L�
�1�4W�t(:k�*La���h\u�T��oߋ|F����[pp6IZ=O��_�|�{�������2R��:_�.P��6�M��G�I�n���lh#+���O:v�n�j#q�ǩV�,�I��������e �j)�D� �i�0(  ���U���X��k���Y�ǭ�3
��� ��V1� ��Y��ba��K�B��^W!�1(	* ח�I�T@���Ů�ks/e�i_Ŧ5��(e�5��A�#t�ȥu�;�;��Lqh�)p��/YS�OSh")�M �B8��!����'�!�C�lXaM0��Q�OgtT���9��V!~��&������~}��AEt�T��%X&��І3J�C��Jft�x���w�٧j���4zI)os|�K޺��:��Sivy�H��4�iE� ����@�)���f�Uw�]今t�
��ܴ�{�p)(Mx���ҋ��f�%[�}�����Ӵ �9*\�*=ȍ="i�5��O����k �o��6��@~�+�M��M����E��������)cK�6�A{��Kp( )����i�]�//C�cV��XZ�"6e�{t�릝�@Ρ��ɋ!�BЅ�u�v�*Z�s�ͼ��C�:y��������7x�V��T�>�[���h$���RBE�1��h��n� �"�nj����ᇖ!��2�4�gZ�F�̦ʥI�6�\����3�L&\jo��
��J:W+L�h��L�����r��G�m=�ംD������r0/!�G�����) -�0KT�����T���}G��V��Y�{�u^��=�p��\#�7]����˺�@�V���e
k���㩄�&�E�L{1SD�4<i�7�y�,�«w0f�z�3���=��#Nya��lYl�3,M�/��4� y�V��-:�2!Xdl� �k��s��_\
�$
�|�*oWTh��]keIᾗ@��9�mÑ�n��[��|@B���q�8-5�>YЦ��<���m��ӨƌH�u]B�lC�4C:��	{�r�8�@���|u�+�5�^�38��Ry����4��3�t�pܥ;���`;ہB���B��
=-oU�q� -4���˙�x����!�%��C�E�a^�Pl�
%�C���W�A��A�� �ɝ ��th�M�Zen��\aR��Jwgm��YT��B��|C���[��a�3
����C%���BkF�r%�(}�2]C�e��|�BDJ�ۻ)������쎸VGPӃU��ƴ*]u�1�t�.~�
f�<���@��FFt:���*��.K�#�����3!A��ȋ:�߈It����j����|��#p�hi�\�k�i]�j�Z*�%�`a�����A�$��u���N�ʵ���b��O�>��꽪�&�\�lS���T��K�{��=ʕ�l�{�IC�g&p�ˤ(Sv`NÐ�kү�Dq��^���'\,T����w����+��j;��Z�%K������%�Ѱ�{x��k�۠�ſ���g�)�|v7h2�1�#�k*�J���]��s_��}�D�MOÉ��{�!��P��R�z�[����?��sf�K�d�: ��8"3�?�V���e��=X���M����i����|���=NBUG$�d�"�UG5>}�g��JLe�Ef�z�[Y6����:"�Ū����½���@����v!Z����X���&�ӻ��|�m���4,��R����J_MԦ�9<C�t����g��5ʌ�	%?��";%s�'GK�Y���2�)���q��ƅ��ڻ�k�R���"Ym6�RzF�
��{�NW/Ln���'���������^�?G�\�U>�*h9��?[�T�C�%����abu��D?����ր�����+�YFG���� |Fi{c�o���Mw�XZ�վ�������l�Hkw���;���*d2H�� �LK��<w5�;w������{�c�U��$��#n�e�����U�����W[��G>�`ͱ����V:t�S����śǵ�����˲�g����+z�����۵J`k�D�-�����gj���d_X&q�!�d-��XM�
wTA�nt �'�9�^�3r��¹l��!��K5iS�D�X�c/�*m��ѭ�@���e�]Y���P��f�5�� +EN.�E��֣����'!8���V��)�M�����ƃ�M��js��柉�M�<��J�d�x'P���7Ú�H!�)-����[�Z��~�������eR�5�����Y6��Oْ�P�T�&<Zi�5Oq���"�z�����i���R�G�NIJ鳨1bh'��24s�6(9/5-
����a�����1��5��g�C�1{xɴ��9a����^����(46�.χO6nE�w��<'���N1�,��,Lm��s�;��ٟ� Qn�EIx�*/&U�Hk7���߲��;Z\�����8��˰���#yg�k�*�V!a�V��
F�z�1��a(I�Uw[i�͔G�+NB<��ގ�M����`����x�.�f�>~\��R��q��h���@!���	��+�Fe����;Ѭ$��d.-<,A.�6-��I�:�O��]h��ABf�ܬ*l(n
z���&&�T�&v~aQ71+�V*�� �;_�0 ��o�$�W�@������n�Bh�M���5���8�#�U�u�S�Ա��.��~�����	�lR�1�9�.��(��,1jߤ�`<=���x���RS~=�Vɸ
��p<n��N��;9/s�2��3�-	r>�-��`���T�ǽ�����N��`�����}�Rp��ge�z�� ݟ�k>���c�/������B{�\�<��� 率�|���9�ƃ Ԣ���C����S�!��...��O?#_��P����Jd��7DD��6���� ��أ���&B|�%�s��pV����M��*2�}��N���4���f��&gn��s;ӓr,�n�p���y�����:9��Z_/ߺ)���� -9�m�h,J��1�x�y�L�'�,�N8{Z0kͷ��Eyʆ���Hg�De���z���q�{9��6����Y5A���m%�hP���b�G�lZ���$�b�/I-O���M�T��~8PUu��e>S��Ĺ���I�Ň)�,���9��ӝa�R0H5�~~�� �6T����u}�~'�s�5��4|M#�Q'�$Ń��G_*�^���o���6�rG�T`b���P���"�,s���.���Y!�.,hf��^�b{���x
�~{��W+&[�׷�|4�Zi�-���6aAEADNKxH�H���#8 "}��2r�A �N=�-ƝM%�1-��]�!�0$
֌��3,]�������Yj��!l�Z��#�`���k<O��:;��D����^֟`_�$��6ow\�E�1�.���9l��c#YO_�A��$@k{I$��A�^ܷdŃ����͊���P��<y��A��������%�줁��<|΃kթ g���$��8�Ž�s�zW$%{7m�NLl�5�]>�P|FI2񹇿�b��a���DYD�
8D�@ a�k��b��;ިL.��z7�ZK�L �������fӥ1U^��qT�QN�(>�(����M�N�E�2��W���c`��ehX���&{ɦ�k}Yr3��7�g�| ��	%�a9Q��UG^���|���	V4#��HU�u&k�D�rRx͎�G�J(0�m��k�_�W�siN��س�	���3hQ;Jbn�c��x;*n��S��<�{&З�� I��G���3Y�ʯ�sw��Xڲ����s=Q֖��O$�"�k|(��g6��Gj�A8�y&g�����]*c��9R�a�"��4��noIƪ��O$J�m��W@O�1טm����6�!xi�R<�>�ř�o�{^RsH�#�H��o�U?ON9 KG�~ds��|�ʮm���X�/���
��|�U�{n"R���i8ȠT�NxМ\�Q�Mc\$�
]��͑��e�����\��E���&�s��}��,�r������y�>��i����w��yZ��x���o.���Fc������ݳ�������@z���h�.G�v'���B֗�"�6�߻cctH� ��ka�ѡ��.���;C��<Ld}����-�Uq4Y^��O�Ǯ�#�K�>�y�b�T\W?����Ęҷ<�E@,����t��[�$Z��z`v\��͈�N�����v� a���]�7�3G�i�����X��U7NI�������PMTp�!Y�t� ��3	��P�~���������,,����xy�p,�M'�������H��B�x��.���*�F)������S=�����)��Sޕ��Â IH\�=��<5\��V�[#r���vH{���p�R ��}(�b���X��4���Rs�vy�_��P�"��a���_L@,4�^�hG1�4��	���Xs�W)t��,'pdW�D;A*��:& F�WЊ�I�g���[.��P,'�w����z�k�j6\�0�6&D�Սϐ3+����P�ZJR�y���$�#�U8��zV����;Tۖ�N��/�NP�i�^��|�J�n��Xi���(�)d��Ƶ������!;�n͋_�-c%�q�I�9L߾"#������pmO+W'��K.2˻�/�^�!�OU� �%�,ͪ����+�m=r+f�bC��·���$B��-.���R�}?9� ?�n\�Ǆ�˅ŉh�qO͍�-�%��^�AG��<�_?�/���0���ǧx��olfK�l���j*�On�ǳi��VG�RR�j�ڦ�nO�}h�:(1T��7����@�3��Ѷ��g�ݎ>�k&����o�!WWY�&�s�:a,T-�q��'y�����>D��̇�^���ǀ
��Y��)_e�Y���Z��_�Q��S�џ�u�p/V����V�?���hY"�3jӡ�w�f?N��)��[��^6���f���k��)�T��{���*��G �_嫪46����M�jSd(�q1y|X��@ƚ�4������^�H�D^�.�{�F9�ı�6����$s��!GI~C��7
?q���Z.ڢ�[I�3;Z��1������lx	�Iܣk������ݩkHCm�V{�d�X�pϱ�ZE1B�{(ʲ*a�R�|A����^z�A�_pn������M�؊�����E(�űx�R�Y�c��?���8b�~�b|rc-ķ���N(��N���!v�4������6P[�%��vb�0�j���C�
��L_;:h�h�Y�#4�dwxRLT�?lU�
H�7Q�ܕ�������AH�p���A�H~jԟ1�����+N�Ya�_�`L�
���k^��('�/x�=hfK�N&t����$�Ŋ���1[	�_�V9ȥ���X�e��h�X�LC�jX5�O<8�=SV��;�C��O�'^�{;�1  f.���V˔P%O��F7���/�����W֙��,GJV�v���$�&�N�jH��gN�r�x�Y`A<6�6WG����o���C�@KvP��%6�G\�SҬX�\���YvW�������l��V�ߕܡVt'�n�>�0��etއ�d�k���p&i�k�ǣWGF�����q�p�b���Y8{�V��֔De�s�a���T�����C��Pڃ�-z��ZzR�&q75�R�蟪Ċc1���hP�[z�j�(䆽\I<�:H
{� -�O���)_���pl���ڛ������
��W���-�P<3l��%�����b*~v#��A^�ǂ���d.�B�?� ?�M�����k��>b�����������9\Áf��c0�X�B�H���%P	��;�
�O*���]Qv8���!�� �I��.#j�>;���	SV�S��x#c�L6�&��_��ؖ{��ظ��WY��ub.V)�4A9�v#;q^��k�(�8B��g�@�be_�z�i�I2��F���{��,?�v�T�ܖF���[��g}0���I4~�y:䭻6 �8�8J�p��c�,�	�bo��Voy��s�	�.w����>�nw�GA@��pV�f�e�F�؊L���3�Οx	'('��*�QfH��.�V��2�rh�C쉬�v�1),��p��(����V��}3eS�4?���ȓF�Ӕ�xOW�ի�K�,���j⩵p$��^щ����[-'����^�$�k	(ӹ�k
[ �S�EBc�!@@�c�����U��Ӗ4y/��Zzx9>�� ?��~;=����O�4<���I`��v�����IO��E��7Z�����͌^c��I\���@� ~�HD�k=]SjMe m�:|�+2#��<�)��s������T!�2c�\i��O�~-0aCb��B�����ȼ��������*K?�>n�θ�O_�<EFU�q�˕Z��􋥡�v�->�%�C0�-�q���]m�8� M?���j�j˖~z���@3,��\�>�?�<5��ܰ��Ꞩ����L������~����Q��%u�Qy�"�ʈ�w`�wt�}��x�Ea���Xw���+Q�n��E�u1���[�{�2 �x(�g�A�P��
��g�2�׋��l�<���F���n�7�n!w ���<+>���}ecD4U�&����GY���0�:Z����+��>��坒��lA*�GC-��Q8��b�G3��7�NV�dd�$[�o���[�9!C�s���N��N��+��hw���⹸�y�Dr2��8yK۫K�����WOT����D&WoVD��w�[�P��L|�}X!^�z̚8���S��qO��jc���>�*��ޞ����#e ��5�'��^�chF�F�8[+͕�%.JHL��m��$`<�O�{��}�y�<��;� ��l����������ǫ>�t�����cZ�է?�o�b�7Td/R�+^�eҚ�Ão��*M��],cw�S�$�[�fCe�������%]�3�܌�z��c�M�b�5Ǐ �캺�vhf�b��i�3H�� �K۵�7CK��3�H��4�he�L;�����.S��@��f�35E��3[�����֔�R��%:c���n��a���&�Go�©���nG�9Q�	���`5	�Ĝ������ك[}|�"����V���2,	�}��7����'5#��e����o;����9�ː~���ϵ����'�#���⭎u����s�a��2bymK�bss�����-A��MN9,L��Rc��vޘ~��p9=�~�HT8	ε���
c[�����%v��5�E�࢟X�8���U7�L���.k��&� �@.pl������D��:+�>��-�ƶ�F�8�;�� ڬ*�f���u^1R�\i;��sa�
U�7���~LZ�r�L�vpY";���b�����뾎��H5�s�]]���,��{�J�֌N+lwr�[P�IA^��C�:��6T�;��������yd��q�Nw3���Y�{(�H�6-�ݷ� �~��n B�0�)U�Cv|Vh^��<q����ER8��.�%�;V�[9;���-q���0�)o�Nt���;e�J� O�C9���J�7 ��ۥ��'���2z[«���H~GC�H��oG$�ee�&}ۇ����!���.Cg6tP�Z� F��c�I&� �a�M��⣠<�fNY`��#�w*}���߂����s�m��e�*4�?y3_�%Kq�N��?2�[BY\�����n��ń�-2��a|\��I����