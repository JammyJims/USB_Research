XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�C����������Q�(���3l�0[�x���l)��P�A�����)�r;F-h�u��\���ba�u�#e:q�-��񆠺n��[6��ʔ�JLZ8�qO *G���j��x��U�墸��v�k���$<섆4g&f�X�T�����y�rM��(C���F���y@��J�*0�7z�[�[W~��]���:=��T��� ѡBF�����?[+���@+�y������2���nE�QFT`��\<��C5
�Ƃ��BJ�_�G���p&\M��P5�)B�gO�@[��9�)�NS�;DA���$@d�9�	 �Od�h=���{�6�2Y�#�,�խS�h�H�nKT�W뤀��h���b#��ߧ%̲:����j�X4��Cf�`����Qw�0�U�hj�Vƴ���ȟ�ԗ�$롣�����['�V ݜ޼�=���`Fw�C(�5�����.�]�sE����Bm�U;<^��xU#x���r4�X���}��6y7TcRQ����wF��^�DW�e��R+<���$�Ł��wL�gS{^��.�4�K�4���	�W��t�{�Z:���	��"��Z��\��>�n}�?��e��A@���o����u#V��������ś!x�|�z�#��Y��F\��t>���C�S�\'W�ݎݫ���Uyg+�����[&���}_P�D��h�G`h�9#�����g@�N��t��h�C�\�%d���z��=�\�x�^}:�؛�cm6w����债kC����#�XlxVHYEB    885b    18f0l�4�:k9x�D���>�ra�8�y�vߦ�s�F��O��.#v�mK���8=6O-EqC��g뽳y��ڊ5q闚��P��Ԋ̲rwl����dO���/4-5_���8lX���c5m�����j˄^#�"����]��7G]�(y�e��:����W'<f;���6$j�v��
����>Ό�\B=y�~��@E�&t�K"鱙���+w�W@�a���S�ejx_i�K�e,�:{t��ƪ�9�/:�f=����4�^!a��珡1�`�}�t&+d�gDqʛlx5r�c���CH�{�L��Q�Ӎ<��D�{�!;�W �X�:+j������B���uvMK���5Q�mc��i:ꍰDw{�Z�����D�#��oi���a�)B֖��o��< ���3C
���rV�G��sKi"��4g�M�<�q��1����@Z���h���W��C�#���n(H!�?��{G�-��]������5\���!76L�w�d��Ͻ�37t*I8[t�)
Q�$��q1�ct�.8%5�=�%%�I�[c �����7���D�O��e�;s��S�R�-#߰BK���{��8]o�ԅQ�~ ~g��y�/$T�'d�T������h<>G�V��U/TQ<:�P~�x��%�H�8;����\��Ԥ�j.d��;0�v�.�R1�������~0�,	��S�t]���y��R�X���!��{ƾ����wus��Y��?�@:���]׳��D�z����)��u��.���	�FLX�ot|� ;�B�HJ��]Q�K�O�8�u���p�>�Y�����+�R^�o�X1����b�@5��S�3�+���X�mn<($pߴ��n���:��*�{�N�
��8/iȥl�=B�WA� F<�t���yr�Y�F2��}s�#U�q'�$Z��d0Iz�7P����}ٶ��%_0�c2��G#�;�&�AJ,}Զ}$�v|Ȧ���	݁ʡ*I~O��){Y6?�=�9�c��X�<��u�/����N����2��)�Eg4���y�d}fGk4|�h�V��;y1O�9�������j�t�q�<=D������ob����S��_��d�ݓ�L��]�r%���xn��n����r1ME���k��t��mvU�y�'D;��r�]�k��y�_b�ꇓ�c���Ԥ�͊�	Gԑ��pU���L��Zhs��k��YA���z�?UwjY�'�r��S�� �姰����`�sV�Lh��7���S��*�#���l����/_�1ju�=@����K	��{��֤��{?����#^�%*km"���(�}�/�ܳ�����d}����?(����`W]��x�Q�dV�}��3OM-��!��r��E���v�ib��,+�y�y�������P�mQ��8���������Щ��f��?�6�fU�f4���)�rX���	��YI�'���dW�aH��o>�#�)��W淰�~J4��3d���������-_k�+��UT[<@EM�,<���m#�ې���	sz��_��F ��� K�n,�KK�b1p�4#r(bg����>`4��m�?��"S>�A�ǳ��7��8���
��,��}���-"�d�%l���Ig�#L=����]p����g`�������w-`Áѹ��g6��p���z�-Ւ&ͻh��>�#|�~L�?��G�*}ѵ�t�!w�B._ۧ��3P��?�id5ܔx���7�𓠄0�+D��f�ev�m;}P$2��G�ėF��YEg�.�zl�}�G#��|T��4l�u1�y�oO}pY����@���k;q�S2X�{/�a��AQ��7�����V ��~�݅�P�J¼��:m]Q~Gf���k�<�/���� �lYU���+�)��gʢ)��1ۑ�o�5�����M��p�m٘ꛋ:�:�-C�U?&6~����E�h��|<�2!px*������3�[�������uR���63������hg�
���.�G��f�5�=A�h<�&'j�E�����������S��Gν����'��É���\ ���`��2�Ȅ�.$q�zM���>���C����^7fX�%��Qj��^;d�2Xmw!���0A��oN��@×�3�ε�d�ڨz9��w=�ș�5�>�p�e��m��xy�ꈄ�P���!�Af�t @e~��%�kcs��k_�v�D�<\m��O��B(f���\ѵ��0���(�⌳J������׍H�~��\�N_�!������ň��!<�2a�?e���!7�j�� !�N�$��7oTE����b��d@��4	*Gf�.Cȝ,��K!s����mc�"��� ���h����{�6�O���/0?s��ee�^r�R�`Ø�a�1�
[��d�F��%x4�8�fZ��N�b�)�8�O���M(�1�K������&�z4B��.��#���^��MNkӠ!^�ɣx�U��8����ůIօ͞Eӵ &g�� ���m��A<6|�ց;o��<_d�
�Pސ��p^��l�@q���bŔ�cN�A���j>K�V-*��
�:!bזh㯂�oVp����.�#'(̃(ьԾID�T'�v��D-��]�l�@�/�@lN�DEDN}6K>;�HJC���(��-&�O��]_?��T��G���5��1���Rȁ]ӌE^�г�Ai��-BB���"{�Gt*���NS�s�A�\�yl0U��
��U�Q�v�Hˢ)�*����bS,)�K2V,B>�@u��oɫB�0��6�6��ؐw1��1��� 6{u?7�z��|ƿ�V��h���'��6U��,���}���� V��!Q�Y�aƯ�¨�g9O����Uޣg^�Oi�|�kaՐ����;5��6T= ��S�I��)X��6�HO�V68WTO!ȫخE���<�_Bj]���W�pj\@Vț8�_0�E	@�8�et���l�vxu�ku�I�p�����U��MN����{��|1�e��=�bI��O�>g�  �B:�T��%!2oTV�̔Va���jUJx�����w6-�U��}�0������3���4�Cg�-��dy|����� ����Rn�>|A�$�7[S7P�o��0��n�-�p�L 2U��1R"Fq�m(�"~7��UX�?�\���4�S�0}��
Z;t��l`uw�Br�S.�Z�ZqÓ.�[x{�}j2�����4���`�=ʇ$	8�D�Cb^U�b�X��3r��$��or�)���{閴�*��A8l� �����~E��*�]J���l�Xv�x�ƘN������}2	a#�l�Һ�>+WՠK{w�h�y7���&�O�!q�A�sl{��H�Q����Z��Q�5,��^z��3#��=�Ȍ!�50�R���p�hEM���F�o' _�7܌���0/�h3���Q	4�|����T���d�2���t�]��m9��i]�uD�U[Xu��aXb3��ª�Z��iTK�)�-��'B���O@��6p=�ݏ�,��:e��}��!�&2��li�1&q��J�������u�F��l�M|���ߜI�Y� �|E��@�����F�H�y�D��>��*�&>g4H� �}n(�U�銮����3��	y A�uՖ˹AAĺ��{��k"�������K�
�
���a��r㈷sA��v�M�6���;�}�t0e�����(���b<�s����~b�.�����	����I�ϖ���4 K�%[�U����6��5��FF�/�(rĻ����/�a�Ӡ�a)�[�)(T�޼����w@Z�~�|g-�#?��	�*zS&��@��e �B)�3J�`PP�Eoh���}o��ѿ!�gV��8��l �.Q��]��ջ m�Zc�-8D����v�7IP.�%c��5�G�ƚ.�}�X��T��1��**���n���aa�(W<T�Xg��j�����â��ت*l^�^r�����i�U���o�p��8i����#ښ�����s5z�Fr/��j��l&<�>KH�l�1p7��]WF�­wcJAW�.��_�$�� 	��,�A���S6�I����F�V=��[A�O�N�a]p�Z/R��W���'�*�����wDnmD�.j�" D.;����e�@3���Ӂ�o��߆������:O�f��_�n=o��fO�bA���짊��$\:��I
΄O=J&iyW�z��3`�Z�����;�w2Qa��%t�(�!��kͦ*���P����mM�.�����0�5��aL�����X]O��s��VD��!(�孇��5��2�[��`�VY��3�����4�]h���CXgt&�bz���v�ϵҮhi9�MZ�~Ǟ�c�ݡ�h�>	����8�%;
<)�܃%��u�q����MeW�kP�j�񧫜-S��#�VK/��MM+�q����E^��5��^�e��?�4�#gȯq�0w��6�Cqw��LH7}�֨}P3��l�i�1�i�Yu��I�+u>6�E�T��uZZd��?%.�t��̧���=���ʍ�n �]�|�T�^��!�m#�1�K���q ����Ҵ���C� R^�<�8�d�X?�aӥ6Xb��DP\cͷ��:� +��|�����D{� )��L���	Pқ�#� J�y��������	[��q��d]�y2k���R���+� :��5��(V,��C!�B�p�j���9n��ͭ�;�,�!�0ia<�8ƅ��n{�lY�ү)(�������Wt���V�6Գ�o�c!��G'�����;��Ac�8.9�^а#
	�����@�3��+��Bt�W��TH���apk�D��d�����Ĉ*	����N�?�j/�V<Y�U��V�Qk��/h$t��UD']���N����S��w	��vN
ڎ!��N�M�>��.�|�=h�Q� �B��Ȱ	j��HwH�NTG��Y�Z05l��/*T�D�g�O�-������W��9���ULU&p�ע��W��g4C@��7K'L�
�^���W���7�-����Z�.iI�vD^����]/���Lh���'4�`�Q������V�q����v�?r�n���4�9	�p��QS4�hſ�C%R�Gh�����_b���������"��Ɓ�T��5�����G�'��뭜 x�Am��d^/������ٓhI�xL�������k�]K�.��O#t�<9�@��2h�t��E%��*�����M����V��������D�A���%�-:�`�ǟN̗�>�(����2�:�dh]�-��C���#}�)��i��|7�����˃X���j�н.ס�9s�����s�$~J
S_�zYCp�}�TI�'t��C�g%�o�de0����}n��F������}n�9��iܤ�s���u-{�X��c0�w7�V��<��+���I�5�J�4q�TZذ�+��S�����3YAuG���ga�M��q�<#���\�ƺ�k�6�߾B��6@a�DF�e���a��g�,h����|1/�����\��wAN�ӆ�ҠY��P��mڎ&�!PFGQV<'h~��^ZA�Ż)@�"���)U���NH|h�N�;�<@��Git��^�}�	b'����T�5�^���R��%����C$�[��Z��-�$����`�$�8��P���~ ���F�G{�R��ݨ�>y���F��#��_��ӻ���������K\�fm\fM�@���=��*t��2�4�܉w�wa�k|��y����VaX	�*`.ܗڬ���?.,��Dyu)�u&a�A��v�(�y �2��������Y�8��u���Z��������l9S�7P�F��xCN�0ݠq�H;�y��#��q�(����h(@ K Q��:�Svj���S'������p�/.��"�i�& MHy'T�����ЎѨC��5�SԿ~���2�k]�囚6zi����80e"� Ad�i;;u���4��
~M����*�w�>��lw�k�?� �o��y��m���?������ d)���u3�xh���n���=�����+j���
ba��'=�P5�^���=�Y|��7Y�lQы4L�cT �Y�j��J"�n�>���-/�Z�n��
�U��Pk�7�Zf����Yv>�FZ��0+܆PK�2�t9��_�u���,ӵtG�Ѻz9bM��y�L_:�TýZ�ma��