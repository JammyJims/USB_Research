XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E�4�^H�va��C�'S�O�_�?��㋳}�,A�LD�������:r�*l�I�pK��l���=��w����!�-ԩ��3$�}�V��'Ro���2�/��W{̑�g���؂�M%
G�J-��Q�)�N���{��&O�_�g��i��Y���VF���e�ׁ���~4q1Xr��1Q�6��W��K��	��Y؊QY�P��4R^K�����E���
n���u���y�^�q4��&�Ku�MTh�6Z��c�f�u	^�'�8�:��/�H
�裒,*�d�$�#Q0l�(���I6�u�y�t����ԅ~U"_��ْEz��!�&s�3W�/��33(,���0W��Y�s���o���T�����*��6�v�<Lb7�k>V����w3����=ճϰR�78�ϛ��V�L���Qo�V��}�x_,�3Q�R���z$}��>#�� +H����/��綁9GmlU�,Ɓ��8=�a~ ܻΩ#��1�ү�n���}O�J����d���/J�}Ft�6ߦ����0Y
~7�m��Z@I''����K@���tʅ7����_�BS���7p3���9�N�MiM��*��;���9}�U��:�b�otT�k����ZB9frL���M�U��;R*��?��"c�/��`W��z����c�LHO:�ș�~0߮���b��ً���{�+*��4�ҵ&��@;�lABQ�t���&z�,�.NX`�-�		�(>jm,s��7�f�-�5	R�XlxVHYEB    d442    2920�����^E����&܉�vp��4y��dopǳQ�:�?�
�HM��D����j�Ŝ���)Q��hh: pU�y[ Rj�VC���`>���+j�8'a�
�'�Z�u ��k/z݇Wگ?��:_YX�z���8���^�6u�tX��99W�]>@�F�l�0W�e�a3Q�.3>��*7q(݀�Iz���v�'��!�e�d7�Rn��q�E�P�k�I
u���g�?���&�]���ɝI��0�=�Cۦ�\�mIꈴ����L�k�}�+�@����&���gu�r�+m�J�V74������ї�;e�ŗ��&7rG��eE��U���Ho4s$F`���ㆾ�A�$F���Y��!#����W1P��ͫ9�\� ��Iĕ&�běc#��r�P^�G���fDj��̜ʐ/te`?���t�&ތa5싮g�?
d�Y�I6�-����4;tCW�s-����b��z@�x���#���.�jf�@���g(vH󃮬�4�ΘyBEu���St�Zv<vǐ�+K]!��K�-�4cwnpW4�̕�#w�W *yZ@ �A�
��΂m����A�5-���UUL������>�?X�xf!�ܰ�,�q��,��.nT��1t���	tT�?�nÃ���(���� &]c�+ �N�ٸ���BW��ƤY��y9��>�Z'ZMh�l�	f���O�K@(�t���"��V�����"��ߨ���ݮ9��O�ʙ	��@(��[4C�
�����ԃ~CL��ϣ�i�]d���v�]�n�%�(�*}��H�w��
�\���'�����"���c3���y�IZ�_?�� ̆h}~�6h� �V��u��N�/ ���t�SE��#��΄֠���
��q"A��(0؜��J��i���T*g���*D_�c�,��Pa��L��t ��=��e��6oi�� �x����Qʱe�>�%��U鼆~�eL.�3�8����I?.�� .�Ħ�A��Tc�9�����L�s���u�����0�g�R�����������?�7xt�Bi�m���i2����j��L@tLSS�W�9)MX�TV~�t+��ɳ����<`r�d{]�Yw%����#XL'�������T���Z�c>Yn��jA���#���6y8y��޴s�x���P8�4 \G��96L��t�i��T���sj�7��#���*�RVlL=�8}c�#>&-&hӍg�s%]�������g ��M�S�Bb)��t8h�ݿCx4��_L���a
��ަzh">(QY�mu覮�������Ѻg���h���D$�-�+iH>5y����'�U�7\��h��{�;oH�_��Dc8j���lT��`�x��VkQ��B���Y�����4���}'>@M�_�=*����k�(3�y^�.��왟"E� 8����~
4n�@%A�d�ď�����l�rJ PZ5���5����&�E���~�	'���	��~{(�%� �N9Z�V���\��,�4X���s����W���^wz�Ί�ܞ	���`x��c.i\K����x���*�?���)f%|4��|��k�� ӎ�)X��%_�R0�Rp�GL�&�1I��u�Reh���.)�@��Ǔ��퉠�����_��<�1Yo�$����e����k(f�4�>'���[�*�����>^o�л��G�n�>��Hθm�1�c=�L��eFi�Y�(f$�b��Qh3g�<���C���7����W�z��:v�5-r�����blV+5@(�`$���^���ð��l�Y՞%4�D)�/%�+^�AHZ��5�P2��x���4]i������7m��N���E�"�8�R�q�����'�Zх"v�,��ྼI�.f��V�Z���Dq"�(%���#��׏��������hn���P�)��GK��zF�c c��Hb�3�]�zfU�x=��md5iB2�q�:5j�D�+0u�W��Q����/9srjS��t�٣���N`���f���^�jJ}����J5��V~��%|<{��s+�D+c�'~�m���ᶰ�j�1�_z�?��D�;~��J������Y��Y�{��
=�1����c�݁~��0��T�{�ی1���=�&*�jMCi@k���67�\1ڑd���m�����,?G�!	A��_Y�"5c����8�q M�ȓ��!���ٟIaw�9����s��@��ݠ�B�)�.��V7�_>M_��&DٱksF~YǍ-�*�/\L����5Q��O�����,��"j��/��M�Z�9�M���jJ8h�qѓ��|2���Α*E��Hc�
&�Up?�qK��n�F��g��g��h ��2�Ʌ��hO��w�grz��*qu�U�_o���09D������� �qE�g��"M.'����}�=}���;)��q0x�U��Y4�<�X>����7�[��GZK7�]"H�|.0�lu~V�c(7�����kB�0S��b��B�/�;�����w.=gg"d��v��xdc�S
7|O�\�'�m(i�tCώRK�ʔ����b_0��c��kS��;6h �RPi�-�d��dYPѰ����;*�$�1N��#�i��/��t���-CD���I�`�	�p�m���Q�,s��;�?�;G��/C��1,��J�H
ft67�gc$���)NM}Hɐ���t��_���SgvH�3|��*�W4r����7<�l�(��F9�Y�)53��_����z��Κ���ڰ�w�{�MW�8S���R�^�f8�6���Jʷ���t;�7�x#�I��)�i.&�@k��Q��ԋ~�V_oǬ�n�ZZ�'ێ�悄Zͩ��3.���$J�a�1@��d9f�17����Vm���÷B��-!������Ҥ{�e������Z�͚.e�[Y�"��k7 Y3��N"�����%zQ�68�ɛ/�'�0ub)�>�
�uڦ���F*��a$ⶦ}�C�Ŗs�o�pu'WAG`�
=��Dc.mo�+�,BA2�zѶ�I�9/lF6@���2�	%J[
|�N���q�"6��5�<�u�$��1"L�����_�VҜt*^V.N#0�Y��۟��;�}���� k���)K�u�T&�虏�<��b��_�;I�@�iV�7��߅
]�}u��ы�S ���<��Z����qJ��RCIVñyM��j�f���1#6O��>Xh�"c�5�����5��7.+����N^l�U@*��@TfE�OI��tHU��ԛ��C���ݛߗ��f#�j6�m��^�%��>�R�&�����L]�^�3�$��p �㏊AC����!p�߫c*{�����}&���'2�z>���9M�p,�W�"�g�y��t����Mz�Y�q�k���_ ���w�!��#�n��my���+]�ܐ��~������~Al�'5Mo��/ �-�I�X�R�>[K�=�$ah2�����3&Ul����� �M]�������)
N�^z���t!�ͩlKFУ	s�^c����m���]rA;p2odS�˄~���8Z������ژ��+�Y/`��h�Ox_i������1K��j*����O��7�՚�|(pOp�|�N��-%��3Qv�HQ�o:�n7�A��C,�B��ǲ�f`D�'�/���ar�Q
�K�_ወ��T* ����L&����D�G!�:khn�1�%�go67��&�փ�n����k����Yն�̬��䦂3%,[f���t��4�aI�0��i��p�i�ǜ�Z��!� ꉃ�B_��-u�g�ˢ�/�Q��Bs�c��`�RdOX�e����l�n�8����O8F1�>?����&~����}&��U=�Kn���<Q��;~7vI:��?}�g��~8�!U�6�B.'$5�"{ �8P5��>���),�9�"o6"ja[E��+�6���)��z^>�8e�N@Ԣ�V�	�6۶B��+�"1d�b�����\Hނ�ޣؕ�0��?��j+���ڛ�!4l�2η]6��WJQK�כ�ܝ� �	�����f�N=q�H^��%Ŷp`�|.�����-*�����B��������pEܥ����D��ݞ�؏T�,��S�}؁�f�ߘh_'�L[LBT3��$5x�(z��@���x�jfG.B��얙�4���*9�Hln��`=
AY�}ש438 
%HF6:Iuvd��.$�dI��.i^���)|�M��β&"(@��M�X����p�J)T�t;q��� �)󾂧K��v9o�;��4C�ّ^mX}��j9 P�=�}��V�1NŜ���#���U%莋p'|�[~��գ�rʣ�a�ؾ��fl�t�N�������DF6<��gHu�L⺝A�t�4�� �bm�BE<9���]�B����y��g����+��+�b��F@����~����0$B�;o݌��#̡��Hd���5�t%:]��`�_K� 洁hV���l%�xtݚ�-T[���:��I�+���͘;}����63�k���u�\�^�k�y�%a��<�s3��Q�ҿ%/���Aկ���0�,���'8�\���9�NLA}�<�c J�q��^��?��it���E�;1�,�;��i�KШ��p+�[�3ؠ�T�9���f辝A����Gv2��;�μ��`	z$���4t%o�qI=���"&��ĂU����!��;��D�P��b�k��P��ש��?ς��[�A�~[��^��".��"����tc���F��L�� �V���1%�C6u�Ado�.�I�<�Y�4���h�tc��d�?��Z!r�fnH{� :k������)���#dB���q���]�ce�Z��bѡ���&ΡVq�/�5e'�k�X�x�������Ž;�C�:��K�Yf��5*D@�<�,������T��Ϳ<�����<�%����\��������ل1'������ϊ?����EK-��fOYEUư�~�?P�i>�#����j�>BkS憩M���^̊��֋r��k�E�'�㙬��}ف]�������_|*ǥi��4q��*�q��t���Mp�d�pZE���^T9��0��#���_�wm_��������Y�o�_Q ���ȞD����  ��ѷKl��"Q2#�p�/ !ѥ3]#��#L{�a���J��2Vxj~@y݀�>����M��<NS�I����I��sX�;��s�ȝv��G�W�CW����5Ol�Y��i@�Z���ka���f^�̔o�� q+_��gc�؂L��`�F㮚�f�/|�eE,��~��WǷU>��]}��{P��//�ہ��p;��NR&��*d���Nh���s�B�K�m*�~�'����e�I~T���3T���G�p��e��֝�q$�)	s�-eΙ|����ӝn��[��h�Wv� �W���}[GK�\�7_�'Tn^ԗ�;T�o�����1�m��\|�E��u����Ć��&1�!S���ݔ�� PS$�MhTU�xs�W��9�}���5&�|��P$�����G W�
D�8݈���pI!����ӂ���#x����}�[���zh1g#��
���y��\|�pgg-�cX�������Qm~� L��L�i�5�	7�d��v���m��eHڴ{��������E�sۛ "���?8���FN
P��n�w�ט����=��T���m�b�?�g!�	�����^�� \7U�&O�ʆw�.�q�%4���-/�kt���r `�V;]輖G�v�;�?/�4!Y�� 58bf�{& +�B�G�����k���y2����4kv��I�nð�o�! ��zʌM�*��0�jj�7!������[�c���V����weX�
.��~��4O�ׁʺC�4�ɠm�����|�֣����{�-�|(�.�0O< �P{_�6U��pDY��P��[�yt��52;� ���
0�*]�K��-�	X��%T���������Bj�$L��G;'7W⊗V)��V#�o�H��j
܌���e��+���w��-z&�����Zw�O���Ĵ;��v�����E�ݙfQ�~ML�{"A�E¯�w"u�Yl�1��r���r�b��z�L�U��!:ag䰞\%hH]�� $�d,?a��ܠ_?�����\B���O̘��pą\(2����s�փ����䍖W�A��U�,��ҝ�����,Ri��	��i��D9iq\�]!,����Eu�M,N���{̩���1A���V�wj�0� �خ
�v�G����j����w[1��U0D�ו;]���!g(� .�	/��|�B��FS��q�U�8e�g)�ٻ��#�d�-S����Zl�
���f�d�K�e�uZh�C����UM���V {�PM�9T%4���@���|�H+���D����4R�x�ނw2���0Q"��XbS�y���zl�ɴ��p>A�2��㶁�,L�0O�ؒ�0��mm�`u��n�t[��M���{y�P�~J5�jin����Zݙ
��#~	��+B��\���>�V�#@io�_��Tv�ӪWqΐ�9��쩡H8���9��FE`��eec$n@T��Q~�ٔ?��%�������B����η�����X#MJ���99yL�֕?�6B2f�nY��c�BC���i�c��P4�h�R2��@=	��HF3_wu�2X���Y�[Z��&]0��q?�Q&�bND�T?u�sKH}o� �Ņ&�א��|r��?ޯm
hj��/|�?-�N{TF���?�ۡ��M<�Ob;�R״�<1�Bf)L=��1j�4يI��|,%�pÈ���e3R�����G�u�3lL�я>�lh��N�(�?�@[�>}�3B$�:Y.����ȠI�1��C�m��V�b�S�C���?l�C�
5�ADu�0�)�AHo��C_�[L-�M�^�R�	5�NR���7�{����HD�����׳�A�o�b��YN��!�*�]L��eՒG��B����F�.s-3*	q�=��В*&��qo|�}^Ys�Y�])�F����z5tg&/X?�S�7�T�(��y��U.��[
R��v��e�h?�=�PS�r#O{�/O_d�����"����LZ6�WTp=�=�,
oO���qRo�����^wvд���j��<̺��* O-����<lG�����rC!, �eBK1�ԇ�1,���[E'C���6�Jt���i��������k'#��^�ۨ�<7}	+(H�r@Hf�7�x�� 2U�Oц`#!{�]'&���f碂9��������=�A ��U5n��)�h����
���1�k���֏�p���=4~ߗ�~�2r����uk��B�bF��O���t�ymf�K)����O$m0��b:��!�y�5�rt\�������_��,P"�����^��[�7��ҥ����o�Jzl��W���$��h:�8��}գ�`Z�e�l뉠�����UHB	'SG��F��j5n$�cD�%���M���X���҂���_SO�*U����i�'S����y��O�t�[]@�#u�/�%>x��'������A(}rFl��I�M'~��܊i?�K�zN��3rv��S��1�:W�C��G�j���ιi\n�~TH��=^����@��~���y�CE4}�F��ޛ�L巼��~~3?����O�H{'��9�ݬLؼ����P��ʪ��fa܌�E Ph��x�d.��	��n�*�v:�
>9�n_�%��Fc�3P{�1�8���~��x֢4!�QTܱ�{;L$�����:�5\�����]���#�R��r4�7*�S�3%�kyc��:H�.��b ��m� ^���֫�0I�kj�BM}���>�4uM}3"��Pv���4'H���i�]Dr��ם�L	T���P����������t��t����ۂ�9aN$F!=}D�g����_�gk=YMΧ�wY��h��U2�q1�-`�?o>� �J�Cɪ�O2M	����]<0�i(
�f��/���|Q���,��@uaq�H:#E�v�>
c�Ӓ'��݆S��;�s��iB�����ԯ����D_��@����C��K�\'@St���r������+�| (،�;:��%$O�'�P�b�wwǇw���6�}�Y˔�R"�P�'9�P�X��"�]U�d�f�m���µ�c�뉅HO%T��'���������Ϝ#H�iȩ�]�p�r��tg)�_)�
�K�M��R:ڻ���*��Q�t>;� ��I�Ǥ���D�#Np��瞜`��U��ay�9�����)y��f�vջ=X�!N�fQ`u��ʀ��H�@�>�b�����R��q�-6�`N���^^�֠�L�`�9"3��������7���2�2�w��󅺲"��#&�m�dX4�5��^�Q��L�T�,��*~tծ�x>�0M�#�j�y�
�l`�l�����}ۋ:.Ie/8�*����L�Ir�ݖ�M���W3pR��KS\���;�+ͳV<���2�d��u��NY���@����'xZQ|�5����i���<$�)��ڶ	�O܄�l&��� A���Ɨ%;��b���qG������+ȏ��,�>S���)�M[^��t���������ξ�f�O��$�6�J�v���l��ɛ���{CT�S��\����&)QN��י6h0���.+;G�J=CF�+��s�/�<�1�8.���ݮ1FV�F����p�j�7���_&�u����}W���$����tV�5���CV}����\��o�����̞�7��^<d���%�"�1)�3v������<( ��Wl�˃���1��)���֡������p#t���8�A�b���ס$�J�FR!F|��
b�La���[TVrq,�5ry��qj��:� u���A.M���^�[lֳ�!-�&ot|�Y,�z�a]�m��=aOV�;]}�+h$�)��:���eNn
w���=�8f�fy�?3��6z�R�T�����֣��N{�.� ja!�>���-N��� R"�:�E�6�R5�#���|�q�ٶ����6;Ow�F줨�:���������މ��	��x��>^%�|�f��A�O�6-A�C,�>OpY'���E�]�9AD�D4�p!UȀ��O�oֈC��>�iVS�\R%�O���m���<���;n&u͚��v����H ��o�3kٛ�@�fH"J�sncMt6t�=Lʏ�j��ف]�t0�MdI
ᖳ�Oh�L�������.Q���\!�[�R�^˦��	&�0s���o$��[�2�@צ	��:�yA9���i������<��=��d��_����R2���`�I�F%N�vͻxn���̇��5����_2��%��<�k[ ��bK�� !b�q[�����߳ҟ	�:B���o�c[���}��[��ػY��FQ㓜!��o�ֱ��=������d@���Bi.�����,K2�4nt�����!�>��~�EV- i�:+�^r7��J2�)��9�!��BC��EүPңHwG������v�sM�ہ�E��V���E���܎"6��v%���~f���n���5�04��p�Ԫ�SD�-�NѨn��q����@G��s���h}]���E�x�y����pk��Mְ@q��`��+*?���
�t�����}bo��\�?1/Q��"#Q��h<}t/��m5_��5��w����*μ�B8�둗��~���5K�]�Wc |e�i�����}f��(s�\��Rn�Q7b�%�	>�r�|�A�~�G�7���Y:�+�7���2����{G�]h�6��1�2�b��&#
��r4&�����i	J�.AaBi�gE����IP��o�'_�e�$FC`�-XP�6)���'�L1f�!]}�Ekؤ�B�]��_bǰݼ�Z�~���i��6�Hr�:�xFO~
�T�0܋~����'�.x
�S��(>*n�-�M�ub�����8���K�J�5���D{�p����i���~<j{~��K/,���P���xeu���M��O�\:�N���lsZX F\��u8i%i����эa�������`Z�^�W�e�Ж�Iw���Y�DLs�1���7�p�������	jn��xA�?�9�^Gq�����s_aW�p5S���oqSp�M��v&��4�U����!U�J��3Z���ү ~���PCV�k�o �����$��:�:2�F�����>8�<���g���?�Gv��L[���c�лw�Аp|^�{�Z��|UJ���>1=�4�T�(