XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����e�Q�GJ��lU��t��Y����/��h�<ܓ*׾�Z*�n�Oj�t��oD�K�����K5o�}�E��M�k6��ϵ^�Buj�5 �T��ME0� TR)���O�����Sη?��7"�9x��z�O0"��S|�4@��.�>X�[%v��W=0ds	 p��c*Ǚ������Ԥxi&8�/On�x}K+���.�|������9�'	jC��Ƥ;,.�tg��'�TZ��?��i���\�)���`��R`*�f@�� �`��:���w�۳�u�[���P-i� ���X�o��<�:5>�zi$6��YߍM'����T�F�[E��qՊ	��U�Ӥ��A�~��n9��B�ֈQ���-���Cq��$�x9�A�I���2��T�XȘ�9	i��bu^��nЮ�E�L�'��z�EWQ��-�e�����t�rّZ��|e�Y=G�0��5�MJr)J{R;?_vc^Y3�Aԅň���k��co����h|����u��������'1� W'n�-?[��W3@���׉�l����ur�S,����y,m[Ӽ^��Y�>>��\S�����awr��a�����<���Iن�k{�B�9��_�&*� ��s(L��fv�Htٳ����Âˬ~�{����:.�"_NB"qW�G��m��ly��<�9E	���F8�ӏ��K Q0���e��v�K��&���<���yׅ'�u���C�5o�+�XlxVHYEB    17be     840��NM�6��认H����?�S#(D��w�ƈ��r< �O:��ۣ�!OE��l+��)K�����F)���i,\��u+�9�)ٴؒ��O��g�7�Iۧ�B(E>8z}�Yd��2F�y��	�Y��3�04������J��6���P)^2��SQ���U�yW�!���K������m9��a��.(YV�yG��íaW�I�q��-�����(��SQ�+l����h9Lׯ���ݣ�/�z�=X�kaA�b�1(���Q�M�楷M]�(���{:��mc(������Y��0�>����_��T`�:x�ьI1��7��P��m�־cH(��k� ��.���]CS����=��|��{�f���
�����QȐ�C�
����D8C&�H�͌��0:"H71�6Q0\g�H?�/%�c�^}��:Y1�����Iq��z]�����SH�ǒW��"K�$�����!��axl�H��X����3��o:� 7]c�T����D�`]���,��]�����;�g�_��0׸w��y`ɠ�[��̞�l���`�Ӱ���{8�3�J-s.zI�/���ޝ&��]�����˂#c�2=��5"`��<�֦*8|�{����R�-sݲ��/z�9�jX�2`��-�D�*?��B�6�&�U Ya��H�L�;�AM�Dζ���w�P��LJ��E=c1sy�͍�R�0ѫ�M���JV�9�O^/��'�_�	]T����DF�"@��'i��2\ӟo����m�0�z��h�q�sNT&����ef�
�Dz�]�#ؕ]�1ɘn��=�H��#��Z���5r�j���D;�/��Y����ޗ���d���q;K�����0�!�_㵶�aU�)@%�Q(�dtS��	��]�B�,f��&�_��'��G�Y:V�x}��H,��?�X<$�w�L���ִ����z\sj'؄�3&V���R	O�F�Χ��
C%\.@���m��P+���˕���~��/�JOO��p]�ʥ�CP?�A��v����YT6�s��_د���<6=�i�<�Y6�HsTe�h�2O
��Qb�m[~��&b�<j[`z��g'�I��r����Ӓ���?�1ލC"��r�a�Gci�O���J>�ͦ7�J��3m��`��ƹ���~+��������t� ���!�eh�p_��	%�Qn�S���\��BL�G���R�òR���T���G��:x`���Y�Wԧ#���q੎����=�2S��^��t#3�+��-�5�f��a�X����9⡦1'�M\شQ�|�b�d_jwwS��K��Q���<����Q}��xF��Vl*�1>Ȟ�߹d�gU�~#�D�Q��p�� �����LC����@9/��(Y���S=}g�D��N�m���-�Tp���];�mm{��{��|�Z"���
;�5�\����g(�b9[�31��{6������5m��/�B�,%;n���"j
hc���V�.F�
�yM��̈́L�Y6�����]�Z��P:���W���:��B�8^���xR�N�J@���V�޶.��T4
���d�)�gSgk���l�����w�X�&��roQS�C=0@����BN�3�]��\6��5F���ͬ?�����M-Է�s2}g?hRm?Ƚ�V�d�v�Fj(��{I�<�S��[ ���Eh�O&?;�qMgp��
���&����pk/���@���}"��wWb��21��Y�	a(�����w��Z�����N��n	���LG7JD
5⌳!mȪ�g�ЬoI%��t��`>v��Md�9�_v�e����f����д�)}cF�ZP��_�J�l7�dF�Q��=C-]�d�km[}�
f�oc�P5����T�XQW�|ąH'�ջ|���4�,�0��%�C ��z*�ONAL ���р��f��Υ�����~�֔�dV ���\:9��N��:��Ps�[�y��8i��ʰ�������Cá���fP���V�����
�{�Hg�LZ�5F���%(C�DE�� ��c���R�