XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��hAL�^F"
0t�Y�g�2�łˉ�+��О�P[C���$y?aJe�-�4� ���m�{���~��ާ��X0�����t�"�Y[�2,,z�*��u5���?�w��@��KT�e J�2����}�!q�BMkx���VU�$�-Lë�(�ZO�`ۓIݡ�$�x*� �����t"D�_ �[٢��1V��z��y�jϸ��n2<��+7 R�G,�>������_+��
c�U;Q?%d�M�����T��{8��,y=+��+�"����'�8���1���X6�[|;�m�ҒA@��֋��,�zAܢs?_b������<o�^�T�T���+:2h^�H1%�^�GJ�R)��+� v���[��ds��ô��s36T۸�\Hؑ��(J3�)KboT�J�QP��X?�n��3h���"o�7�>Mk��]�m�� ����S�K��P��i�n�ܤv�B��}c\�?cɜ��;8�~�G=�����gn��S|�&R֥Q��, 5�w�+T��E*��m3lW�Vb�B���'���u�Г�eY�Ά��*���R����d_�&Y�i2�h��U�Vjɋz2t&ꥁ�X�j�o&Z?�#�L�$v���;R1n�c_R���� ��M��b��ѡ����@Fn�[;p��#Yu��4�	�.�u-�#���YN�L��'�Rܙ�%�����t&��8�6����^{z<��J�F!v	@$-!�z �˵��G�lfў���wXlxVHYEB    3970     fe01s�ޡ�jc�,�T�fs��@!�v�{C
�����>�|S\!2�ռ08���j	��C��V�}�|
����omX���[�BMQ��렡����@ܟ�}���K����	��_��4��v�Gסd >�W�,�r5i��Σ��9�)��K���w�"3x��G0���P2�ΐ17��?N��ŉ�������i5R���L`�_�Dz��R��D�%��v���,X�Ho�/�EWXO3��:t��Q\*n��W��GE�/`&�����(kkL�o%�w�4#��吜V����
��<��YG������`����Kv��u ���4��}���w�SFA	����J4��A/࠯�a�����|�����;�m�ףW<��Xl�I��1,������N8F&8`55�C��[[T�{v�&Y�t*��҆��=�i�漋��%��Ů����EF��IEm�~�� X��Ӥg@SI�}�����/f9�o��2o^0{�����yR��R��p6Oչ�m^�nSZ�<&�=��+\b�=/�s�x��.�[;�؋�%o|��=Rӊ��p�D�p�HAJp���[]�-{�����o�U���d��%���^K"���dYn_�6_@�>�ƃ�bd�G,��-<�lFO诏j�����N�=�[x�yFa����j���4��="\�!d�����ԭPz�5n�qۅO�2fê�#n�3�<��b�>�׆T"spw�I�$�����4��������U�e�q<�
x�1=]���Z�  ���@u�.6��I�����_m������ᅄ�/�up��P�)������ph�M�B{9 ٘7W��o���69	�*�/�{{F���>]�I �c?�p9(���߉O�C,��ߔC�nc�/vy�DREq} �J,k�,�>�=��\��O<c�fgo9@�m���"����ؿBt���n`lȨ���ʿ����_�����e1����tK<�(>��a��L����U�CgOh��L6�e�lI���^g<16u�l�]�"71GV����םA��1��ٽ�M�l�ؿS�#�ɐ&���^�9~y}t'�%�>$!�A�Ռ� ���p��L>G�mޢ�C�e�=`!�X��01Q*o��w��� ���u��Z���NP�����Do�W6#գ�_�5 �����,e�q�澻Zx9+
N�B�q7���q�0JQB�|+��Q+�p㴀�6�	`��%��J�?�w��h2��~ﵵ��	 j��
(
F1�D�U�Ђ�GR����1�S	��ޥ �Cv�'U.e��C�xlcF��]�g5}�.!I��B�&:�ܰi�|!<�������%�U ��a4g�� �[�f�ź�A-� h]&;ݑF����*5��u%<2���qz~Ո8mj<Ư�p}�
�"�5y�	o���|��S^+;��j�����x��z�ʹ�,����C�R�l( >���o�G22�f�*�M�Y�7��%�v4�2��`n�xo��X(ic�w5����6}���}��vq;*ji��!ʈ����uZ�t������!m:/K���Q0lU�U�;t�޼�5U؛R���'����w����Q�s�q�-�@�*#s��{\0�H>����H�=g"���7��ug��4�[ �w����
M��h2���'�%��V��P�Le�v�V�Zd����ѱQ9L'��ibH�W���޷�ްU��T�@�(�V/�JA��gg?E-�n:*�D���e-��2�;��.��B�Y�����&jST0_��T �#���vx+�cg{~�(�M<��2�� ���:�	@��m������z��������#��+ܛ�E	�;���[��Ƴ�|���x~�g�3MAxo�hE�̫�h�Z���e�J�%�y�5�j_������\�׎C�v�@|��ڼ��D�sY? u�ڊu���)���6��s,�g��BW�!@����͟/D9�_��k�CK�_�5(���n���-�Q�]�{���3�\5؅��"������l{�)��+�9vϏL�k�S�Zs�@�R�H��U2,��Ex���7O�
=a�*��{��j�̙��H��(�)&h�@�0�����ϓ��/w����.d�`E��4�B���߰\���y*���d��2���}��[��o�1�����l��������ԚT,�g�����~�F��訔�6��R3�����1����2D�M����>�T�yt����'g���6oa�p�"&5`�'�g\?J��j���`Q�?E�X(�}T�����q@ޡ�:��\@�G����U�M�M�Q���Th�j���8�N��B�(��p�D�%4χ�1Z�m�jޛ�>�H8yzep�'��G�"*������U�ڤ����CƔ ����/h`kM���'#�.Wھ�}�|�.����DV��=(L_�ɛ�Ґ����@�FN��>tȖ3_���v������-s�h��&:�}��fF0_��0��5
i
zj��c��9���P��vc�ބyi�p�i�#���(ia=%�';p���7$Hvf쿁�v��j-�g�=9���9qH���@���fz���XN�¿�����4!���Lg�����l5���"m�g��?[��8���J(3@��H��sLF���m����w�kb�3�����-�X��|:��Q�^=��o��M� ������d�x�����nmt%��Vi�3'�DH��23x7��׭Ѩ��^
7?���㡴72o?
x8�ͱQ}����ѫ�b3�����@98r���:�9�e���*�
���c'�E�XY���'�L+;�%���eu�z����,Y�����v~^�G��i<%�R�����qxj	�S�4J�F�@s�bSE��#�'�9_������3	���W�n�����	�#�y�
!F��tQ�'l��t�_Ek,�;�'^�q�뇨k��`
9+%v;ǚ��-?u���&}_�1Ǿ���()*Z}_�Q�(cY!��.�R�`I<����=��kw:aޯ�AQ��A���78�%��$f���h��Xi��( }|u�fP�c�K�į <�%�Y^6ތ��$P�)�D�����{��$)ur��>��7�;���ޗ�>E�斍0��?5�<$�L`i�S� $w�?Y�~�s�8)m��u,��J�0q0�Os��*����6f}�w��
�q�P�ղ0��+�u�8ǯ1�v��b�3�}b�#\��*[��P��)����ǰb� ���]֟?=h��]�!�"&������aI8n���4e�y�:�� ���^EZ!�
�ʿ�����l�q�D#�R^��&\) ����/�sM6�_����@����k�{*��8����({g��A����_�t�v�.q��{�%��a��.A�E�#\J5���͊-T�0�_�-�0��y�#��}�Lfl)b�[��vC���/R��Z�?�	�a�������dw��}��$Wݷ��:����h�{(y����)���06X��\����jxj�'�߶?\����N
���)�c擎�c�y�o��! �	@pJ���[�b�}�]T�������fC�}�
kόo�����OZY���I�W���{֫V\ht
�� xj�<e)�;D���;Z|ɝ�Aڢ�����5�H���WHޫ������%� n��٤.l4'5�*�֦CheϢ����'r��!���9z�R�o���_���Na����tr���lu�q;B�<sچ�+��d�v�
��v$���i�L��)8*R�Y�B'D���^5�

R;'> �U&f���n/��<�U���RI5����X{$���gp�Ɏ���PTŰn�*U��m� ����F,�sb�����O��~����D��zr�p������`yUz�>�ogy$t�=�
e�D�(������)}�54��F��,�Su+a��ڽAy$�lFI+`yс�