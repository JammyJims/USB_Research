XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���׳:O3p�sN�K��8H+�꺆u�McV��qȷ���*xf,�Rn��~�$b�K����rs�j@J̒��_i�����ũ�%lJ"0>��F`;�V]��%d%O����Kg)t�RLV���&�Q�~��x�X 1�#ƌ�,x#���O�r���:��>���=�1����!g��s�:�ێ�[_#�&�u2�[�5�f����0�:�T�)P:b�K�_�ml�|�G�>�{8Z�l<:�0�;�'$a	v��D-���	���W�-ڤ�F��T�};��Gη8��H�����胏�����(�2�Q\��������
E~�=s��.�"�P���ȎL�+��	�&w1⚳���e��H���W�D�sC�=ɻ��>S"�7c�@H"
�m��N�p=!��k7]��1's��y?�.<W��i�����T0�ݤ��
AB&�t�1H��`�?�g�'�E�� ��s��aB=��p�[�F��1C"��0b�ԩ�@C�^��l��_���R>q�%p`ʫ����is	�oY���r�AK	' ���P�P����,k^]^����:�Bp��/�Ay���1C��aYj8ٯl�T���q�H%�
��:�x��U�R�r��_�F��Oq��^�S}�^`�E��Z>o��1�/�q$�����6Wo.���3�J��4�z��/��,S��O��kf7�V�M�"G�>�ӛ�mؗDq����.CW�]�	h��z�+t`���tc.����XlxVHYEB    20d4     b00�N�oc������@�p���(�ٲ3F/�<^|__�?����Q	��!�%�����U�ϖ�a����/y]jW�wsl򦦊-��9���.H�gC����s,�y�6u�k!��Rz01>���>�1o�>W'_��p9���
����G��	KXt��+Z��G�|6	���x�=�w��zSxɘQ*2-��v�1�V]\,��g��	��r���gNYa�<>��'�a��/����k|u�leL�>�J�@�B����UC�vm4��d�w+ZJ�E�9Wd����+�N�/��z�{ܷ�I�o�}���+{�> )�Ќ"�@0AK�C̨��r	��(s��m^������v���a�ϫkڿ��_���>�P�"_�I��Z ��/�'�f~��5R�q�K���"an�EG+�K�vJ�"⣢S�3m&UK��_~"8TVg�������%�^�'<��ˈ�u�����+���(2Q��+�zo��+P"��^0q����@���8UP����@�s��������yֿ�kx�� �)��`��ܥϟt�4��+����k���B��	֑���~q�Hf�h�8�CB^5�q}�w�6��u�_�R��fVL4`�R^�1�\��Ŀ��g��9�N	��\.���#�|m��-7#/��aF��8�Ac؉-�,��6i_�FN�?C[.�� +n����j�]�����V Ҫ��2���[g�P΅�Fb:E����wbH�++�L.U�Q5�c��O{��o���m�TA��F4��3R��"3�'o�R�>^�� �Q)�S��+R�>��J7�[Ց�5@	����#��g�/N�i���sd���M�1���yPFlO��8Nm�6���^��d�`��]0k�����|'L\LJ@�5Õ(2`۞�6�����N�iM��k蜕���J_���Q��/������Q�.�DE�H§�j;��vLOrӹ�������C�!�nNm/�o���Hb�V
9s %X�Y�F�2ò���G���FTū��-�m��Q�~�{*�8\,�̐7۾A�%3�R+���[E �ֳ�ë9��h�\����x�����=�<�l�8�������x�:u�����w�1�z;���<����Ϻ[��5z�H`�)�ݻ�D��k�O=q���� W1K�����}���iq������P�}&�Ks�-�2�\�@���x�n|��'kT�^�Ǭ�@Hv�!յ4'w�q�28F��|C�Xʆ�����6`��7(2U���fP��%��~��u�<K^?���[CT�qV6Ǽ?���z��W���l�Q#k�8~2	����=%a���KQ=�^��5�h�
�ZkL/�?�RL ���F��v�sQ��J��0uF%��Ju�7�JM�V�T��G�n؇0=�^E���M���8yY)�i~;���`�p����w��[����2�#��o��H�+�A	���LI&�8�cX���a��?�����"q��r��?<�pt怇�0σ75�g�}���ېѸ���H�[�P�<i�~X6�L6��>]�`�5|z�L��\?O��&̃+{h��1�l���h�R��U���N!�9�{�Q*U�E�򦺦��u�����f����y��VE6��Y+T���[����7U�mB��$/q;�G>Y���C"��y��&G�|:�r6�)H�Q��_��M�oz���pPu�YͰ)�rʠ�=���y���o�^B�H��A�|���.S��wPG���JL�8������J�{��Ę�2'0�)	�8�������Й �oǱ�?������Z��8�����z;7Z���[j��2#�3���tAZ]Ňb0�R%�o�ɨ:2�D����ӡ{0�dl>�7$Izm�����vt�M����N� ��T�L	��"6X:�r�A���YHV�����_p�}�y��W�!5�o����X���RU�y:����c54a���+��r4��B��ڮ5�����iDVfB�=�(� �&&UY��ݛ���F�9�j��Y��@��� �x���Ƀ�y�>;��d����,��S�PF�d%��	��ob�U�tZ.�X��z��/��z)J7;�B�0�������.��׹emPg7�C���N"}�S37[�J˾�U��B�ʰ}1+���N�rc���k#��x���q��/vE�-N��&���e?�aDM=�J�k�أ�n9�h�[z餐f� 	�Ϟ���f~`8~��x�N�2gF?��:\&k4���N���N�!����L-��m�6�.����"�&��t[�e�����ߞѾ�~��90$�'����6l��ꡁ�|�ɤ�7�d;z
��ݍ�?))2��>���J��u���U���s.xo!�dy7r�2s�x7�G���(�����a4Ƕ�Ƀ�-3KȩB�k�P(�t���i��.�7㰹���3�Ќ��c���Lc<b7��ał�����������;��w(�S-aπ��S�ݐ���g�u.v��ߩ<�B��$ѩ�V&	v[��i��p#��Kc�^"�W/Z��2�L����`�z���,�= �4��Z��:�5�3r7.�S�_��f��ݑ�>��W��Ԭū3�"�Kj�a�j��ڦ�(��I���\tht����s��D��^gS\��sh�`/57��g8-���i&�|H�n1;n�Y��&"�9)"že���#���Jv��,�&bDn�V�2��\B�u���