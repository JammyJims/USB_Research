XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ӭ�U,���0&��M`�s�s'g��'�0ˤzv~�x��͘Y�2���y7�$Imx@�X7�{-Q~>���dX)%�sF�֛�ϫ�:�����_ �z�+����>SGV1"ϯ��	��~��z���)ۃjSE��W�
!�w��E[���������D��Xu;��5ݪ\I��fS:��Ð��0J���N���d1����=Z!..Oށ��Jxe:`e���5=��Xp���я��:�f�aAY��^�e��4j�!B�q;4��O�}��wsp�[�2u��2���$R�pbME���+owVvс�Sk"OnPV�� ��\���_�;���E�}�E�������`�uy�����<7�	����@h.�sW�\����Q���������f���F�(���Ь���A���&/5�O���Q�����L�M��X�{ҷ���"'1�~�qd���E�gϻ���gگ�n�~^y����ߺ�Tݘ����֟s�|�z��8ق�r���nw���î�H�53�:Up���Rl˙��M��
$ޝ;�^�g����4g��kv�^�J��}�z ����xv�ީ>o:7�\~����G��p�r�Kb��c�����%Ap�ί�Y�L��f�Q��i�ӂ���u�Y��S���/}f�]�#4Ҍ�����V��eD�i�{���EyX��t�!
 ���nD}l���T�5"��[�h�Y�S]`��'�fa�U��t�l�XlxVHYEB    2bb4     e00�\+������;cv<�����/JPߛ�jB���R��oجWx��|q�����^�������vv*�^ɍ��wٔ�Ѵف�9�N=���e�J�����a�w<{�Mz��ή�J`���Q�h���ݐ�bM�L"NY���x�q�����UA^46̣6��h9�E�3xBJگ{ʹX��%����	�"��r�=Z�mmO�wՆ��Bm㺄`�ױ��aq������K
�햆L�_��<������%��9�	�P��`ZF���5�pr �
$�[�<KW�e�3m�6{�c~�ھӳd�v�/��X%甏>"��r�R�k�
��#t ��)�CS��<�K�^��4qƛ�$�,�9�J`G����l@���4����b�'+ �\?U�=6)%�,ؒQ-)��8r��5�gyz���:�(�i��A\������<�S๪.s�=2=�y��T|�=	�Gԁ�u�K�����[� a$�5���
~�>����N�$$�%F�<%9����ȡ��l��͹�蒎���N֑8�3��R� '���KM0����-�/׋
ߖ��q7�*(���5��.� I,l���sd/en	�Wa.����g��Kf�Z}�D@������#����[{?����Ѧe�$�M��<m�fӸ�~�4��-_��
��!�%��g0����oZ�!ʚl�<̆`��ov6M]�9}�@�_kh�{N�k�~,E|�
	�"br��$�v6D��ٻ�A�B+�:�Լ��^�z�,�N}q{����p�0*�IӉ�r����Zw�)2�.�[�o}|�����4�\G�������� ����7��kn����!F�%l�N�*�$S�BT���^�{{w��Qi��:��X�
ݽ��VXd+�&���n�L�)$}o������qw_�#���l��̊�Rl�4�d������{%�kR��	V��%i~�/���2u��!X5�����c�=^�/��l�6����9��E(��v�YUZ����|
Pv퐎��!i+A�� ���1�2�2��D�`f�^_=���^��k���55���E���&#��%�;@��#$�b;( ��7�c8�ӊ����	�?�)x6VA�s��50�ц�:���n,�7���N\�D��.�s�2�U��t{��+�i_%Ĥw�sj��}H�ӏ�{ep���?�2	��7%_�"��L�ݷa���+4�F�����6Pp������(Xo&hˡj���5���%��V�(e�Fpryi��\UBG(�<��f�����"g�,7�|p���cSA�}�}�
��b.5����1˼�*Q!���*���sv�2�n�vBJb"@���k�M��f��⧈��3��09��D��� !���5A���p�%q�d~E �"_�R��ϯnk��}6���"�G�҈'�]�]�Y�q4¨��aIU�ݛ���P�߃p)�iC��bzB�)%���A�<�N�m�@Tqp+���s)/�V����A@<im�z'�ױ���:�Rg�@3��+u[)w�m�,Y���<���.����vN��}\l����V=�:���r��M�@��*�j����I�9�f5i���e���D1��z��,HZ�	�]Y7)q3�ן��4��̓�{xю�l��[L6� ��RP�å�q��em�R3�iX�I2���<Ja6��D���ML�ݺ|ӕFG�Gʁj�?C+�\�OOE^x5 7�	C@$B�1oe)�2��?���ֶ;M6ƥ��&��q���rR�?��S���L��)V(Þ@R"�����R���u���v�Ե��Po#�gM�␎^:G�?)�����7z�a 1�V��k
�I���*�ӱ���c��e�ם%��p�i��o4�ZT����T:��𕒎�H%��C�g3������c>X3D&�f+����K��F� �4�S�1}���H�3!����*:B�kd>b��V[�):�ȘC��DjU��]��5��;K���Sn��-US�g�΁@z�B�7*�a`r�����;�O��^ �8�o�����z\�#]�<�1�<�.I�-�ܯ�\���3H�K�fE� �:���x�ͨ֟q��0��(��Ě�%�y>���T�T�yY�b��wQ�c���F����tA4"NL��w1�i���S�,$���;�~' (O0�����q'�����oUY��=��p�x��3^W��	ǹ�V,�SV=lA�d�k'_�2Dt&���Z��%�Y�����*�H�4�����,��pgs�Jw�υ�9>]*�L��|�=[Kw[�sԛlZGձ�|6#�K����0!��R�h���8YA[��X�0:	e����>�U7��)�t >��]ľC������֎��M���ϳ�Xo�U���6��bG9��$��)��MqI÷�����Y���6Qs�P�] ���ݿ�u�?Y�����b�}�7zX�T9���J�Z�=��n@�\#����,K�׃dC|�������/n]G�������f�T���P�Cޗ�~�
<��/��ղ!
����@��[�������a"{;��i�5~���m؟w��'�o�+��z'�o�"9����{N沔g�}��W��x��1����fu>��R��<+��dnAa!J]��F`�ʑjT��zB],�$�J�w�W� w7�N�*@-E
��UDׄ�t�����,j�~��ӭ�/��&��a7J-�S��v^?$�.gU|�'��^&Ǯ�Ӕ�LԻ����u�2ȓ��d�ě�M�O�im=��1�{c����i��>؍`
�wb4�Q?;a��W2�*��:q Qq��^#�z�Du�]ʽE�5>��&2���na?�H�μ�P�"n�^��a.��BѠ m��h�D�.� )�H����fk�i��qm�"��ߕ�w!)�Ԕ�<�nS�~��8r��N=7�ey�j��]O�N�2�Kٮ�AZ��G#����G2m�U�=�~m0ϛ�v�u��V���3�=m��A�C�m�zy��������Քc������x�C]d�y�8�$N4U�NAK8�r�3Ɵ���V�������G��=�dل��Q,�xW�n^�,�-�򯪍UT�RFՋ�ʳC�@g;GM���d��T��9w3SGYc��èK��1	1)�®h?S��A��0fZ�����$�ǡ��5:�$��Tw�8��g������Ệ�k�t+'+�Up�{`�PTu�,��	�����j��6��I�4� ����Ҳ
s{M�m�a�gd�A���4{��tg�*�2vd�A���y��$\&�`�,r�������W ��T�2"���~�?��y�����k�#ej�)����\��i�#G�������m%"����.	���?��'�`A��|��_��W=��i��#����s�t9Q&�ہuA��~J+AV�m��|�|`��M[#�dW�e3��J�{��a�x�ǘ ��1�5�E��G������̟�^y�l�k>����� C�ae����"��'-0[