XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��uޡ�/�G���:k�ܡ02tn\J������(���������5ZЇ+OW:>�]s�\�c ٟN}��K����WBJ��cq+ߺ-�#�tX��D���~!�P\>�iB������ɝqb����1������z�H�����|V���[5���F'�$�}BtsI�v�wx��D��` 6+�GM�,������8����,��xnf�����۰���Y��3�/���;��{5�t�=��Kp����֞-`P7b�Z��}p9.!s���F�f]B�a��`�5|���@îj�����"�3�ӝ�7�T��O�k�U^D�I���x���;� H
����P�p~��هU� ���>��2�$��&�ʴ��������+S�.R�������T)���r-��\7�S���� ���1��bW���6�����70�c�9�`��Fu�	^�����){�^U/��=��,��j�/��ۨT����gV���G�����^R�"nN�#⅒�'UƜ���ͤ�(�ɠs&m��4��g�� }�E-_��j����|���"�f�쉠��5��`_F��#�:ʶ�-;5,����aL�ʻ3`�fr"_>�^�$f�ˏed��r7X�E��v��0o�1��A�
�R\X�0>O�M
�Y�V�%_ƅ�U�o������Ɉ	����d�?(VqSf�02(��տZx7X�
B��Pi �rK{�r�M���ٯ��5�������&$霄%XlxVHYEB    12c3     7c0')+�B��ĭK\k���MC�T��43|��.B�VD)8�g]?�a���F]c*��t��.e���휻1����;'ň�;�cm�y�ٙ����T��#fs���+!#bs!�8���_���cl�/1R�Z|ǣ�y�	�xz��
-����$XI��me�{����#g�c��jU.�����O��H��}�D�V�k[���vK�7&TV�g�P�:��Uz�'с�f��E�f��N�9@�?s���o^u�~F;q�e�ʁ�������AQ�-�Avim9X�!3��d|��C6��s��[e��τV����J�ڼ!P�BL�����z�9@ƻ�(���o�y�~r�9
������KB�b���~J�o�Tmе����$�p���a�*�����(��.��0J��������������'wWB�_�� rB�Qt�XO��=��.o�h����m�]#�z0�GK�k+�"�a�t�v��9X=�t9�����%`tiI����y���G:�G��s8pS�.��B!� �/�m!v��p��:�BS�4]��М�y_:�Ї0�L*O�T��|`�EM/tk�[���=���r2]��������JݎM��q�n�4-�օ��a�~w����F�c���$t��s�%�N\�\��9D�h6�K�V9	&D���gw)�(>(���3�t�/������D;���y�ܯ~�K��Ӟ��gW�CPߒ�*�L�~����P���&@>޹g���;�����腣sCg�&��3��m�R�jߩ���gQU�h�*���R�Z�.��Dc��uÿ?L�7+���<�+|�5&l�2� �8G�����8����C��W�;/M�
uB�����0��F.*@l�F!x�@�;�QQY@�L9�Ir�Pr$�ŧ�â�Ug�n�Y�WJ�;��&d���zi;���	#~��)#5��Y�L�G5)^��qwN�@��Dw;�<�F�}�@��U�{33�.0�K���!I��u�%C�]_ �ȉ�7$�77���8t�/����B����B}jw�V5���wq�vFt׀�A	B�k&E�9�0b^��h4��\��Q0�
�l�~��k��r{�:"}�?f-���o���n�]o���[��ON`uݢ��s�a.�s�J�7`��oB/p�I��H��7���m�&o��*\V�|!l7�E�!]mmZO��NƿXS~Š^6z�~����2�B
Cȼ�6�/o�M��c���]����Y�O����h�(S'vXR?�K�$Zf������Ѻw�����5;�Y� �KŢy^����K���[�6>�vɈ���� E��lm�����Q�b�Х�ʻ��\���5�~q[ o�	�ԺuJ�H
pi]��-b�1��(^F���92��z��D�����x�G�9`��Nse�VG���h����]���;T�Fl��� ?M6�Kp���15xZ�d��J���t��J �� �o�biֆ2�kz����d�^U��'�Lt��&��i��%��(��(��_E-���5�?i��Tp_ug4�6�X��h�ֱ�a����33��2�#х6c��H�艼9_��IjȬ6�sv�~E�?!9sjf�(�F�vٱz��8�z"��Q}�qs3[C i����t4G9^N�~}���%
����ߙ4Q�m�Ȅ�7Ű���)��z�i�q��D�h���a.xO�g����=���(l�� 
���`z0kT�e�'|�g]R���R���Y?M�|��mx*u�4up$�pt*���sa�ΊЕ�z�&so�y:M��e�?T+䃧~�2~AA����CA ���ÙP4|U��eh�u���KL��q����,|u�aD����i�!'������9�F���+g ���߮L��}��:;Ύ(�CӴ��) CX��[;���`�����}�����Q�u�z�Y`;�t'�J�g�z��rT�