XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=V!�!��u�����_(I��?W3:���k4Ğ���~�؁e$Le��p�F��s� �[�{~�n��e<��ܸg�p��z����xJ�a��$dQ��	����*-,�=�w#�܀��:
d��"�t@�2{j8L(�l}�Mď�,ddߞ���;������-�S]��]�־��A�]�l,�v6Dr�ҡ˚2H��������=zmGȘ1aL�?�O�9�c`!�:�x�����F|��������M��р�s#��"	�躹(�6�df�T�L���aC���p`�Ku���"��:�*@�S8�-nP�M�`���"w�"ju��q]&Tm.v;J�t���X>e�Ju�G%�Y=�S��7��I��@���c¨���k�M�Q��!@������<ު����wY�6����\���"���+]"f�m��J=Q�o<?�+a�ƴ����M����ۆ\�=ШP�щ�Ȏ5��~�h����}�Zǟ#�k������Zq���̔��SRݐbTq�NsB|	a�EG�� ?F7'r$�u�P_�k�:y"�@_p"�x�C���&�.��B�I��d9�-{�w�h��0�?ۂمT��<'nR��� �Ρ�I33��/S�a����GL!��/�Y�k#ԕs�:�h޿��)�=���y��o~ҥW/�cow'!BX��.�7����	t��ـ
�����HÏ���p�C��P��]A�UR�c�[�2��\�Q�������L�U0}�Z,U��AXlxVHYEB    144f     840";Iŏ�oӢ��ٹ��HTx��J��B��O���������X��q_�<�d]?��JM�����`F�g�f��{����&�\:�g#�e?�TVB�¡Z	��1�w3�4�ѧ5�����w�5�G�ܕ?~��ki�p��;5�4�����z(�:����&}u�d..,�j9�<�E�$�B�ׇ���I�;��E��+��b��؄�d���H�˲�7����@2��6���B�9�1�	79�^8�Oev1M��<Q�N��{	,a����E|<��!�iD�<���"�6����^�+���*'b�O�_��7����j��JS�ڲ�]8� i�~b����QKg�υ��u��Z�Y��˦�$5z�Sې� �t����X�>���}6��0ۀ6>g�h���^5�$qY:
�R��&�3�A05�,D����S�l�đ�U���L"��U@������A!X(��+����Ƌ�'��<Kh������n����#���~�D�T �PH�S��*�SĜ�[�	 ���pד��l�3յ�9��K�@U׾�)|�t݋M������y)�!2�J]!O� 9l! 1�o
L)��Ϟ�j]�	�����u�߿S�Ϗ\��]\�����0G�9����V8�ټ>n�vO��]| m�N	�S����_��,���Ps�U����م���e�F+�� X(���7�Q�=��!˨���%&���wv�.�.�����1�KHq��!U�c��C��M!���3��(�C�i�[�:���7��\��KLl���N�s]����B�f?�Y�����A���T�rũ�~��N�[����2�2>�����?�q�q��d��-�qa=����^dk����S�`pm-\�%�:t��y3��k.u?�k]W�kå��m�O��=��P��NTM'{L��^1��~1UjG�wO9A&�EZ�ceU�Oc?pL�B�O򌲳�>>�I��˪���=]�L2��Y|�j�ސo=y�RR�k��L�W����&��6���8DGJ�P��z�34`:�(�(2Z��U�Ŝ��6w��I�H�@�C.ob�2@��?|�5S�����! P��ӥ8Ċs�ٻ�dL:�� �{~Y�,$@&��)��z��J"�vQ�Z�����^:C��3�?�&/�dD����@i�?:1��,��z7o ��8�1xZ��48׃�� �����|��%-�:�<S�ņ���㪰����H��+��uΚ��mt]�[z��4�xa��� ��H9��	��_k���l�����|�~+W�^|"�W�d[��T��*��A�a�|>���h�}w�9�V9����ˌ֡���
��Jl5)}�!���4U� ��"h"4
�&pg���9�b���jg�~'~��)8h��\?Uv�#���2S��\@�7$��%�c��K�������V^�7��UV���[�jn�69#���ޥg|�$�N��/��Lae:�myΫ`�rR=ږ�=�|��n�k�i�h�6�j���<��y�E|��Z��1��>8��NH`Q�"o\ӹ�x����bq��������*�A��X%C �avX��[�?�v��Čq�7��t��Ċ�\=�׺v�g~0�"�=��R�uk�k`�!>�ֶ#rt�jm�� �g����"{w�>ܒE������)��l�Y_	�۱���@�J�F^�0�e-e!��#F��P�~��&�7�ۢ�f�W�yQM����	]X�y�s{爲|��05�58ĝ��yn��L����b� ���,\9��1�{vݽ���	���9�`{�w�7�Z\���r�'��D�!)�;z�J����o=-�������b!��`~+h�C5�9��=b*��f��J�c������@~b�H�q�x���^;��y$1�\�\���n����vEj��	yNھ���%�ݞqd�9ۢ�!��כ�U�+����3TS�'�xML�E���Þ'����P!�{�p��+:,�F��,���L2�T�O�f\�.�G�f76�����H�����~_�k��8��Ţ<kS�
�VlU���w��*X*��