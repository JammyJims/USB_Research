XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.�� i2��.@ݷ'b��Qc��a}�U���A�c������t�,<�g�/���4S$�]0ٰ�;֋�6��.��
~�H�0�F�QՁ�O懑���#�`��֗|	�X}�t-�i��ms��O��Iq&�%LO��KƬ'2���!�����0�-�@�_�e�;=����n�(bV���X��J�FOB4����g����^���^/�����0vq�-d�S�����<5��\���g1ځ�:Ӷ�9�oz�W�~e�k�c�����ɣ��x�R��¬ۧ��Dܽ{�)W�E��u��9D�4��>ux����R��)K��~��h#/��<��`�"�E�+�`��h����)���a��R����%Q0,Z�m��t.�DY_&譔�~>c�PO��ȪT�[3�*1"+�eY-�����h���;V��>a/��(�?ݔ2�
����J��/c�5�����t�.�&�]�-BaJ����0��M⒱��q׋7�Po�E�!�B�_��&sks+}gD�Tk�GQ8��u����L��}M�w�ˉ�MY��"J���֞��F��44kC�!�����@�@�+�@��9|(��$o�0xE��<պ�C
ux�@�> ��Tm��PX����	/���G	��E�w)K�G~�p��zO1=���z������������}��g�ڣ��_�;}<�f�W�=�����{{N�SFq�Z\e������_R?qd����N�($�(�=2�lk�^9���:4"�A�XlxVHYEB    26a1     ce0���S�ﱐK�U��7�%��T�ο���)>�2�{';_R��ZE&��/�?2@�i���EÈƦc����	;%�U���z��'~Cn)����	( 8�l�֢ͤ۫V�?Q��(�Ί�CX��pq���Wq�G-,WŖk��pSt(*Es��Ti2cc��sS��&j%�9D���m�7�#0 t�H�XV;�$�R���Xk]����e<��}�gj]���(�J�"56Ҝ$��a�aƜ���3���Ҵ�� ��\^ܘ"��@Y�p�[��1���m=t�U�@��HJ���l�YL���9�����e�P"Cx��j�kh:7�-�`��0{�/��{G�+���}a��c�f!y���=�h$S,�߭�ɔ%����n7������7��:	���M�֖�Ε�$��7qpf�f�n!l�����@��r���NƩ��/�J�(S�GŸWs�.?�O;Lޢm~�(a����n�A4Wck}S&TF����l��+�&��yK����q��:��|/K;���hX?�Ԯ���=�,5A�7�ޚ���l��/Q��#�g��|���*/c�)����%��èO����
T�>���n�p��J-F���x�"?�ԗ̈́�r��m�q	P��G;p����Ү�:�c!��2O�6�+�g^:\�d��6� B����a�Or[�����h��*�a����11o�����l��������c��G3Ϗz�i;��W���_r�bQm90��p���J^�����/.{�a�RB_&�^��[��P�+�*�K��h�y7�O�ƷȜ ��g�]+5��)�*V�/�d��Y�/���F��1o,PG�4�AE�=Mh����r��b� S��Wƃ:�x1P�Af�sL~��ۀ�����VН,a7�\�|�[}��%2�wU�V:"ۏD���M�U����PY�7+?��z�$UT��|����!e���8�B� JW̿ y���Q �I�E��&w�������aY�y-�C�6P(����1�Jw>�A7-�K!��`�
L����'!ק�-[0-g�M��=������vCβs3����#���O&5��ӓ�F�fԹ�V$U�3�z������7&k��+�?���n���.,��+��e8q"��S�
�-^!�̰>��RP3��3{Qp�Ea�nX����|�����lsخCM&u��)-�|VΎ
�Ô&y)[NB����a�F:4��p���TF w����Ť�$Ǉ���U��ڍA�E�AȑLXU%���F	>��W��A��D����i�()�3�!����ҡM��T�U!���Rpߡ�����ϩ��K}�x��ȃ붰]��_ީ*�8M���I������&~7��KØG����9����k�4��p;�Mr�OeRy�r���*�'$X�4��bŉ�ix�N����4e�0H��K�����+���=Ē�uc�B��x�/��I>��8���F�y�k�iL�ۮ�*�ά�A.A�6���2��ɣ��O���7�V�d�#5K�d�5k�,��PCy��WP4�z~@C��<��٢Yb7k�����[�2 �I� ��/%�k����!5��c�Б��,��pa={�|Ʋ�i4�0�&��$�o���c���@8�E��7^�:����ZO�3K<�A��y���Zդ�b�b��W�
�&^�1x�c�����
�S������SmriI	�L�	yg��|)�&�p6�x��4�
���{�yu���5���Wx��)����~Y�Yb:z�>�2��5a�FķG�E�hZ�sf�.��%
l=�"�J]���BsyQP��m욑��h��W��[鱽�)��,Nd/؉��h��=Լ��Nk2bI)<�m�@��Am��U��z�G��.���N�=����F@��$�?W�9m!�k�0�瑿8N��t�NO�X����º��h)-�P�"��?J�b��ғ+���>�����S�l���5VJ.��$�(�����m�j�^e6�I��|r����?$Ӷ�)Ӏe�qR�:�~�y.�ɚ+�}�%�,�iy�&����^��4�7�04<-�^���7E#�ަ�� �A�lo��c}�	=�%!
�M��(7q"QVgu�D��y�B����=;��Q����N�DS����@�`b��G:8��;b���F|�r�ʈ1ȖX���tcg��[�,�2GA��]M_nM��E�K���t�(Nj���L��D�����1����/s{�N]�-�S}C@�N�	2�"����y��[�hD19���P�I�	H�Y@�w�;R�E����(�k��`��!����#D�1H��7T�\1ţZ�MK��tы���6�p��@@6_�ۤ�N��n����h��ep�&��d��t[��L{_�{�"��D��[��.�R�Xoj�'y)Y�*	s���4y�K�W�de_n�r���7���U��������GĶ���R�V��`b4�C�����u���.>��j֤Dǰx�K�k�ߢ��fK[t<��R�E�ۮ ��cPT�Q���{��[��D�K	v�b- J�T��䲔=<Mn���\צ�1���{��W>���S��f|޾D���s�,u�p�LЈ�y�n*�Wb PB��ag	j�$�(���5JN�pw�=\�Mh���:��~���Q�<�)E�|6[�w=�U�����=�I��V��-g�4p���6�( _��b��u̜��e����5d��Ր�?%j�0��N�D=A �F�o�]��J�a\�� AF��\p����9�bI�R�wV]�22bkA�Є3��(T�R�8�cj\���	�A�J�%������Ys�cʷ'��L�C��v��tJ3zR�`��9L�?�4������S�;�`��v��N�Yqw�><�m�aFnm՞��i���C��M��U�;{�2ͦ���{�������A8E�Y�R�,C Y�����@׆��iS�mFH*j5�3T���Ov���Ka��"�!Fl��w.����t �D�*���4�b��Ŭ|E�Emt�p�+o'?�b���l��w�d����e^pN� mCG4n65
�G�k�	�R�z;[rw��J �x�%(�*�����$�|�w�%�Ώ�Wvz/��%�i�[=%�T�s�X�Sq6��=��G�a������s�����Ӷ������L�?���p�OHLMqҋչ���s[E$�l�T��