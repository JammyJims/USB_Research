XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��.��m��ֽȗ��6�;�鬒�>'��<e���LPO�2>k+Ԫ�4T��#�Ee+���׈dۏ��IK���0Ń�5���Qo�c$���]�Zy���"bW��?'�i�:Pk��6� Y	�(,��ۙ�6q�>���l�)�nH���X�р��	F-��,�:�k�j���m��D�gQx��y�q�
�̊.�ޢ��-�P�H��^H�s��h��`��R	-�+�T/�}�`�nQ�>� Ҏjↄ�9�陝����7�L�0�C�N<����s��Ռ���h�%Y�e[������@*�|q�O���y�.�fcv' A���e"68�¨��Y��ISZ�nԌBW*5f�� ��,��?�:�����=d�	���V�\�Bױlr����C}��=x���?�by�S[��-I����;�f�CMԾ���Xk��&�h=�g�w����q���˞.&5Vw�e�υy� 1A�o�E���,���3����`�i1�mL�ɼ��zLH�Y����|Z��9݀��|l��\̈���)�VN�9�p[j*�MM�syO������W�uT55��t�H�!�H��ڝsҳ��ʽ= �Zλ/�5�U��+t2RS�Ƕ��W�edٍB��x ��ub~��,��!�2�E#%1��/w� M��"�_��@��83�IG�����1[�qjböv��`�gO������ii�sf�v���z3J� ��7�eԥ7XlxVHYEB    3282    1010����?A9	~?,sjLI`�Ta�w`�t9��q����=�.>g��'���YF`VF^㒨;�������OX�!�g"����eL�-����/�v���C8��BgX���)�� =��<:���qI�a}�]�����%$��%��#�WP�0�J@�ɦz>����wo��ꉍ��y�K�Q��WH���ut���S���7��՗^��i@��}����O�(|!+D ���V�;�i!�J���R����i�d��`���|�_��'o`�eR��-
_H[�b�4 L��j�sBhXX�Ų��ͤp~�w���LY(�կrȁ%"��?�L�)UY�E��p�-K-���v�UM�_�*X��<��V�vG�6�2s�v�h�ڤh�%��H�xʵ�\V�$�y��L`�ؽ � Y��S���xax�@nNw�Ʒ�уw���{�
ʾ���ņ�fN��׸��3������+5�H�ߴ��h`�[�y<Z��{��ç�:y��Xv�X�^t�O�g��n�~�
2���<D�m:=�^�8�!�_E�2%��yᵄ���]~�PڑE�S�\[|Y������uc�7|�In�Bɐt��#���Wq�؈I|(&�`j	h�Һt.$۶��#�2�Gc7�z�A������rm���{����,t2�N,�.��__�lr��X��LEh��H�v?�h�@�i����A��\�o�q�U��B@��ð�n��]�_�6U?�{���]	674#Ĥ���X�Cw���+-u����˖;�-ֲyr�	"�ZḠF��9��?�w�?B�{���{�G�S��������ꤙR�Ƕ�_�)�4�9�����~j����##�z�^�Տ*u^b�P�'�#�T=+"�2�f����{�ѫ��q���&"2�,J��Z�f�����dks�2�[�V.�����X��3�`�@�ԌHA�/H��v�X9jK�Y��	��܄G=hc���90f�q��j��rw'2���������L�%*�"���NW>�]֯�W�8�����g����B�NSշ;8k�8�b����J����
_�<�]�NH�W+ί�����6��'+A3%]��c�#�&+'����g�^�
NFqN��S�'�V�35K���P�y9����R�n*�(c�fj�JL��WV�}Z����nZ2��':σ�_=⏡�L��o��h���� .>�>O,<V���OEb_ϐ0��H�?h��k�Y���<B�Z<��:����
�w���,D��^+���5�0�ʓ��˥�Nw�z��IX@��>1?����w�x��k�Ῑ0*wkEl�w,l��^p)���.B���)*ZW�F�w�3Cn~(\մ�����"4�ԯ���1������!�%���EtZ ��a>�A��%�s��ef	6��!Q�O�r���9��W9�f4$lL�h��>��fſK��XM�Uׅ�+)��k��g��:��w���@�Ķ�\�CVDj}tyI9BV՞�A��O.���D
�.]�ߡe��&�.�<K~Տ�X(�4$^�G���]��m�� z�:��.�m��rs�TS�o������5�7�T�x����$�ѹ��Q�O�~�wbAli�5P8�n��#œ��GME�֍��s��n�#����a<������֋��h齱�"�K��g/��q�'D����
?�|%�==��\ИD;"��cp��-�����6�1V������rQ�Y����$j�0Gn�=f,"�� �$ԳJ��g���7���J��X�k��a�76TMc��OЪ�i�EE�$%`���=N�þ�xV�)���������"_2�LTu5y�e?^����'=��P�%���R���3G�ef�$+���	%��V!�'�Y���|�������Zs�n僝<���{):����qd?�E�o2^H���N��h�����<blѬ��m.�$q��S�URm���"�2{���y>����Q��F�6��û+s˒E��e���h�jЂ��2@�I��9�1�u�r��D��g���ۣ���`���WG7�",�h��N(�48�����k�"��K�mzȚ��jm5O�RF��kDf� A��g�X4{�,%���z��ҥ-��:��@�oQ���C�-��	heM�-S;����:iDg	&Hn������劘������u��V��>�ړ��;���+�+��G��q�D�G�*k}ϝZ乖D��q
n甒J��A(y}X��S�R�:8م�7k]�-P��Yݿ�Nv�ݳ�U���,��RvD_��8�7)���N���U�M\��Њ���^�z2�������O��X"pٸ�S����ņB״nz��e��9l�J��鿸�1�ӑ���X��\6�x���wMn�2p@�FǢ�*\�%�gl9q{e����ED@5 X�RDF��2{�?vPyI��F3��3Ⱦ1L��E���T����Фh,x��M�)���������vQ5����`��77[]�_>l6!UN�^9�^���O��a��Q�
գ��2�*�����V���2Mm���Zɿ��`5�#�-�'`�%|���^I��Ԕ.����]C�⒪�ĞfS�sc��\2⩆�KK�G�=+\�Ȧˍ���l*�b?'��g��_$1%��������C��,��(�������f3f+�mw�ȖF�8O�T��`g�R_Q�I�g=zނ4�eaH������eŢ8��w�b	�������YKY�`@�)�N(ϭӅ���D�c-A�s��, ��-�~���EQ	da���y�h�6!����1�#�)�����k���u�t%�z�z�����L}n�e����=�O+XA�C�5E�Y'�I{�z�~M}��A� Q6/���.\�S6�?��q��W!>�>L�����RF�k��J��|e�ٗ��Maܤy�TT�|�'��g���c��N�g}��Xچ?Zeu�ԞXQG!뿥�q,g�ZTر��i�%���s��0y&T;�'��/�9�0�N��%�O�,������ ���+��MR�@[�;�Ň-��
r^cQ߇�2R�O_AHaD�����Y$��@f��2��Dy0Ӳ�)�6��ᜒ��˭%�G�.cu9�Q�r��4�Ȗ�( :����P�q����XK[�a�����8{2��Nn'�j�Hy����!�o`v�qf)/+�t�&������������{u�.)8�OE��8Fe����>���&^��b, �|��;�u�6�GV��F�sGH�J+6���-�����fƍ�RңY1�H�#:u�C�����W�.".�ͳ,�M��з�s�ڢ�������vk�"����Mb2٨$X�w�u�\�J�~��~bc�v�v;c|�����4yOCn�\�rwX�@{U �s���WeR��Ui򬓦P(�֐�S����
���<����Dc��9��}�V>������W��tC�'4x~Y�F5B���{��س5��RI���Nv��yj�0A*#!����:�E���H����LK�������??,l�2��0Ձ�Y3��W�!BNMd���5�Zdr�C�B�*��?=iE�D�S%5]sF{��T6�9Rj5�P�W��
W��
ϋY=���o9��҄#��
̇�q�=��9(��?����zy~\�J��mc5��b�H:S��z�C�㙍!�|Q�cB&m���fԂ�	��V��_{3oCE�١�T0�e�O����E�W~�#�������]�Y�E;�-�S�����w|J��b=�<���n��7"q"^��/4�#È3ί1���	,)�,�~��F�O��Ҙ(�}dN\�A*�@�2�m�'Ykj�?�ӗ��]�,���S�^�Pw��O�1��Yh�K[�E�[�!j�߭�n�geD����[D�F�W��\�9�᥽#ӗ�?��b�I�w�n�"*	�h�)��lb}=�Ό.j�8�w�
�D������X4[��{����]K4�bO��P*�F�X�&�	