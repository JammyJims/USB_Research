XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���u,ߛ�;��N�Y����~�
�r�K�GW �VC�7�|���w�MGɴ򎉖=z'�M� ����vf�vL'8G?�EB���]���opj~7
��J@w�|����v'�����*��	����x�u�ɺ�E�_2g�u�Yg�;��F���m�fO"�pV!Ԅiӳlg�8�V���:ǣG�Q3I^s�-�p��T��jC�N��Sq�u+:��H���kOy��+�6���T5g��Q9S�	�g,3����+etӳ3hj	�7`U��m۲���O&s�����)����́��ɞ���D�T
��⹓��NEUH����+�~-&��r����7o_~Y�3�-��\5f�i<�N�� ��C�Cϋ����U#���B�5g|���"y�d�6�U��D=�bNB���~��VC%��ʅl�
-S��w�pŝ���s]�ɵ�f>��ܕ��w���vƉ��*�8�x��͔�ƊM-��A��|�f'�j+{�Y����Y��[��@c{�~f)|7۞{؞]�r����^o�NF���^��:�S��ʸT������j��mӅ^�\��ň�7�4"{��ㆽ~���dV��A��P�?4G;vn�=\x��h�����c��E~x�%ˍ��D��c��	f��	 ��y|��W���Ԡ94I�ױIk �K��l㽭�D�5����5y���÷���6:��ף��
"'!I��5G=^���W�|M�Г�Ip\�2�U�'�G��XlxVHYEB    193e     a20��n����� ��$��"eً�\�U���1�j[q�/����S�$VGm���"~����u��<h��A��2��@�]织G�!S��Y�.��KP�H���:�y�,��/T-�+�dW~S�����߈R�p`&��5������P�X;q#	d��˪�SW��Քa�5���kW��5|%���ڟ> Y�;�8����9�~cM�Q��t�V�v�[bi榥S��t�U�ä���4 �}��7��(A����n6�wg�QB��L�a>嗨0D(Q;�3��P�W� ��^8Y1� ����y�S7�����$%Xz�+�z��y췿я1���0�[P�9IL��!X����$��L'
�J��ps6���'�|��/��K��#4yo�wWP�%O�0�.���R?�M���B-'Oo_%��w��]&��Y���$�����z2�OM�g#ā|���J_|*����)bP��{���b.!٩��Yo	/�g����p���%sC8BЮ{�\��%��gw�ބ��Fn�d�a��KƟ~u�rO퓳CZ��v�c!1|�L6��)�S��f�l}~�zp�?n����H]�!J���ј���e��؟?}Y�
��asrĤ����I��r��*���,�ְk�Ha�����8�Zֿ���+�������d�y��i���Ğ����|���A��MG�S��vg�(D�x>Q��&�Hi���X_���8�������Aq�����aE8�Kq��?6�y'�%�����#n���C���?�:f���������ܪ�C�8M5��߮)_��9�xI�����؁+UK���%���Upr7�p?��'������?��u��	@x(r�3k15}Z�ݰ?i��I��������b�^I���0 ��S�Q�oS�B�.Y�i�J��4�?%?%�:����(�i7���P��z�Ԫ3�Ԇr�������$�S��v��p�
*�U/;��� z���T�rm�$a[��j�}Kk�-��ah��>P%[	z9Lq�1Iߝ��_���@ْ�/lN�Y��],� �$Z1�C�e�3�%���E��O?�$V�Y6���B͠*�h�`�c1�fQfG!۬���w���~�X&	���� z�
�(�1�7W������@rߑJ���~�ǽI�V��`������`*��j�[�nM+�nĊ8�q�f�1��jW3ŝ\�ꤵwd�t9���-��"�ܕ���)f}M�M���)��=~�E���7ݶ����j�<��6�4�Y���p�e������{��X�����no��a4z�BJ���'tU�V�w�s`E(l� v��C���+ܹ��!* �c�"��nJ����eؖeu�k��h2�W��|BL>|��o-��Z�Β�SP�d���o9���t����ו{m�b;�56��-
���������bAȌ�?���"�}��w��o�Ot!K�i���Z6��XD_�ز������\v1s�(�+�#rQ��+��S1,H�u�ĝ�+��SK�i918g/K84r؊B�BUI^U9���EY��7�9�9��z��X,8��*~�)�JYxu:�_�v�Z�����H��x�	uRt.�1��lg��ڌ�$�ff�Zٷ9�+dn�[a����Ɩ̝��Al/{�i�Z�F��w��~Q4��R��E�jh�,a��ݓ;$��4�2�A1�|F3b�P^@jۦfRpB[f�}�*��"D�����~Jel8O��~�D���!�Tj����SX��vC,��c��ȟ]
mb��u#`���?�UȽx�Y9^�}A����)�1&�� Jۡ�	��5�%����b�.#�7�Y�\vj�E[��q�nN�S,�ɯ8���eM��I���g���V*?m#N�J�Fց����YMU��Qu��K�H�ۼ� S\��ϖ��yظ�};0kY��d�3*~д-�I	|��vZP��(��1#6G0rvM�ܔEkkĀ�����ZGb���{���R&6/DN�Z��p	��i�i8�O�r���c��R��Yك`,[N�dU=Z��G5`��>m�	���K7vh��9_�MU��i B='��2m�G��,)���@��(�ˏ��W)�i��[�\p �.$ɓ?0����~̔��5�D�=���t���j��5(o���!7+v���䝬޾J>�6q�F�R՝�v$
�l��)g��`�@!�T���Ms%�7�A*|��S3'YO�ti���nE��f~7��.O��Z��Nac?�ؠ��u���"���$��ۍ̅�}������,�[JUq�G��o�e@�k�|MJ��iiU���������(|��\f,m3�e��A]��
_��gqU^>���K*R#�]�.@şoW���2Su�:�n�n�]ߐ��4	 XP[�c�-V�S�Ȗs<B`+� =�ޥ�c�� v8�د�����|��f�[�<,V����Ӝ��b���<_B%�~�< ���e�y��w���߈�z�n���d����0�悍?�'�.��_�s�Zn@�r��l�l��}��G.=�\�qF