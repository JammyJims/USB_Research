XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9�^��B�H��]�X��މr{B��<x׸���f��G�7`�>���n�/[���±�x�#�o3"����S�G�pG_�}�������̗!��P�߀tz��T��,��� �)3J�&���hYo.��ү�c+G��;mdF�:��S7�*=jq�(D�vgضZS.f�j"綋3gM$�N�#(�s��	��z�:?���j=�XL!ډi��T�Q �O�wz��o�+�j�����|~C�[R��Y)�f,	8yC��uLw<�����bТ]�)=��D�h��cOO0?=YwpݬϪ0ꢳ5Mm�YH�>E�H�l�p� ����
?)��Y9k_�Ҥff&�:ԃ|ɝ�ŀ1ץ�|i�����UC�o̢]O �Z>�S�|�3�Bl*��5k�T�������S4�o��5(�?E���fTjx`��	B��3�*��/�]-R.ۓ��q�����I"��BɁ��V��1Q[*۬M �#u?0��b��N@(m�1�7BZ���bǰ�bզ�%P}�Yrd$*��4�\C�b3:�[7W��S�5�i���B(i<v�6D�Gu(��-�z��l�e��#x,3�d^$^���C  rS��9�P~QĐ�ɏn)6�
2{^�s��d������j�(7˙�Urs�]��MZ��:�w_��qrN�Ձ�2�^ Sum�|}�ex�50�]~� ���4�BCm�Ʌ���QJ"!�����hW�ZE&��y�1`���{XlxVHYEB    1314     7f0I��9��ҫ���:���2Vhf�i�M�u���\.'�ceGmٽ*:E]U�NÃ+VLnCQI�v�|�Mp����ME����?�<�_�HC<<r����������<�<�N�#��(��'��V�l��KbҌ�A�pv	�Sbm{g��Ҟ�Q�u:�����H~?��Xԃ*���	��X���%�7���J �'���f{�3�_JHn���o<�_B����0N���[b%�֙M4�˗kW�l ��M�ù'�a����{ď���@R;�I�l�!'������j��3���W��/�}�i5�R���/'��gw<���|4 ����!��J��>@v�+�1ql f|�~�%���C��Z���ܗ2PN��_8׷�����)4�)���y�I��UO�it�d���D�r��>��(ޜ_��n�"gҡ0A �Nb+XV�]=;�)u'���s�ī+gs7��DI>�'N0kq>zڇ�H!���ZQ�`"A��+(�8_v3�o:��i��L��ZR?O�:�QVء��Z{�
��!-2�~}�Ӿ#.�
pUt�.B��ǪPT��6|D&���������}z���}���_�].���ǐ�^��+׺�o��n��Z\�|�*s��O��	��D. ҇.�-g_ ��p����x�K��͟�~�7s#_Xe�1����J����g���������R�7&�P.�]�S)g��̪�e�"��9������7�b1�XT,�,���K%�*'N�k��-�p��/ �7G�F���<{ɷ�K7܃N�u�0 ��R�̯\;��fc*�\ҕ԰N#x�N�H���������k0�����d���3l�^�2�/�[�A�O�Y^����c�׵����iᰳ���NhL#gs��λְv������ �,��:`AE��- �x� 5���HdkEP��*=�s���C\�W�ɾ,�L���4����Y}�Q�*}��Iq1hw��/w�Q`}#�[	W�(�����+99*��R��'
8�5�Zf&)�7]}���:��A#�h ^�@怒B����iUB���(������OEt��M�g8b��M6p{m%�$�E�os/�������K�M@sb"��b�Ὥ)nk`�����`�CU����6b?��:4�i�� 7��r����q�*���^���OC��^�
3	���<�W�4�t�;r����^������@����0�0�JˑH�.D�W�f�"Tf�7����M������mCC%GyMeǿ��q�U�y6�l��k�ϝ_]����K��1RkĂԿ%m8����ǚ]���lM�Z0�i�4�F�N���Ax����Q�|���Ԓ~(M^R4����p����M{f��D���^f܀J�"�vP����|��d�c�����������G�?"���R�j�6�*�ˏ!���rҺG�_�����~���q�@ݹ�:5�G�*�%I4��J�{��'�ƶ��)���.s�]���ނ-�!�[�����;�k�L���)I3mHȺ�îv!�~�N4�����:��a���X#��/�[�m���.D���w=؆M�Y:�sŦ��1I����כ���ڕ
�p� ���3>Nz�bD�C�7:�QH��z��A����6�s}X+�*�ɣr�fN֕�f�^�.�Ěf�=�1Ǝ]���[�bt�,X]��DůC�ɉr�P	O$gr_�QJ�k��^���g��/e��A2�(^a�JR�ã�t�$-eo
'���$�\���ܽ-m���R3_,���M�����Qe��U4���rF�j���E���������`t��>�]A�����lX���;!��@�
�d�f��.R�S�tO���{�OG������v�AO���4q��sL��s��Q5 }3�t*,�ѰNcS���P����`uԇ�!`���@ �;B������5�#�Gԯ!;���ӭ4��>w�ZB��<���7UJ~;x�&��X3��`�k��0P��