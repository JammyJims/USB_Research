XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�nU��8��Y���ӵ�	�4R4oY&��zi>��7\B	W�G{-߆<k��&���@�+mӪ"aD#L��Y(,D]��'瓨��U�_5oR�b�(���C^B��Ф�u5w�ą�ƪo:H�dZKuRS�0a#�4��r8n6F{��\uTшJ�0�.��S+��#��yFǖ}�!~]�l�� ?!��M�	��Dx��3����J�cJ���� ��h `xD���]8���h	��)6hK�?m�H.@�u�?�:q�s�<��F���������RUۉ9�/�IB��Z���ϵ�v��D�dU���2[\�8�'~.u�vհ̟/��x�~`���B 6Q%�g��+�_^:�n���T[Ѓ�~��p������1��LOO8��^� '�CJ��!�&�b�_�Y�_QYՉ"r���5/R]5��:�܉���1 1_�Ŧ�f��9�A�D_�z�G�W3�{��0fS.&���P0A�rq�q��-
�s�o<�,PP�����I1�*�9����bWj6�=^�����=��7��a���*�ڤ�y�V�1���v>��B��/�&Myq���e�/��bZsx)6�[:�Z	�c��8ֹ4���0��g�
E�gf)��i��-����;�Ӓ8�r e7uB?,���dp-D���X�����t�0M�9�����?��G���×��T5�vBJ�0��?��҇J��W_6�V�a���.�O*K�n�c`���
K�_���W`���s�􅺵Q�XlxVHYEB     8a2     290�|����Y��雒K穹΍Di[nR�pH;�ܝ]:�8l:O>�?$�kf0�{;u�q��F����|Mb���i_�xk@zo*lڰ+9W,�C�荪��'4aK�'��e#�:�T��lvs��Ro�̵����?`�KtC����<ѣ8|/�:1؜�Vɮr!I���Ul,�%��3bY���3���}�NM.�|X� �� 4��e�N5H�E��>�ٞ�EƓ�j�|a0�M�k��1�@cH�l3���L�抚��PH\��>�r��Oc��Gc��@W?��
|�O4��O���_ g�x�ʮ�ǚ�M�+#K�L"���y�&XU*pG��S9&d��ϐ��H�w���h[�d&�ϧU�"=w�6� �������K��*/)-ldx>��A[�M
��=���!��:���	3����c�g�`
��	JP��q�iMT�Ƙ{J�u�D�,�r�� @��'³�"1__<��;�h��ֲ�el�[2/6�AZ��2���O;%J����M�;��b���V���Dӑ�Qvp��Zb~c�S+���/��#�w=�Pi�>e���s14�qb��ʨ�B�7�lާ}��X�#�(��t�A�� v/ƿ�B
;y_�-�!2m�X�W�����MاG��#��ƌ���/�V"bav��E{���&