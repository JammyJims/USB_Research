XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�6�NS�K��!ƏR�#B	j�U]/b�������]��)rߜ����ͻ-g;~3����ZG��6���{�9j�l��o�=��Dc~)�_��J�9����= \�[r�)f'��-�3$�_a������8y��3YO�F����jb�3����F�@|(õL��w���5p�yN�<��@e�r��MK�"��,���ok0d�6�L��0��*���ۃ�]���)�9�y[�_�{O��a�Z�|w�#�W��B�:�w�kW�%H2e�L�^;h�{9�bF'�xO�Z�/�`ˇ��Ŏt���\�l$tq4��ԟ-�N�_[�mf�����8Y���8�t�4�Ɲ��F�w|sr��4셞��!�	����pfWg���GI���r`і��t-fXPv�E�O�/e��x��5����/��*�As ��iX���ؠ��&][�+��)�eB�J�@��{bG�Y�Q��"��a>k�Ha�������E[�v����]�+B��?*�!�}�a�4]��ȣ�z�qu�����$�>sW{�jv�T$iuĸu /��%5�L#5k���
|��ӑ�4�ȕ�t��  �/}<�U~�"��/hX+�wfR�FϴLA��9Q�W~i���� i�V3W�����߷x�sU�a�X!C�����B���b �3���Y�@��]�Rϓ��4��k'�"|�X��>s��><���� ��CɁ�ks�꒔�̒�4�l��zW0�UDXlxVHYEB    4a43     ce0���?\��&������M�v�V�������<�ӝSn��������7o!�]���#�h?����=^�BY\���&,W3��$� �OpĜ�5.!ԙ�D�&�m��N#}��<�\}�O��� I��$�_��ҙk ^�H����D�S��<,.����9�3I�%���"���[01�Z-t�	tVqO{�����W�M)L�B����*j�k����$vn�n�R��	p4�u�$ϕ:��˥%q����K��3�iDs����Y���@Pcd� ���\�i�:��?j�k4*}��knC��L� ����jT-[|Q#�£��qc�v�L|�
�D��n�Y��/��[lWB�!~��(�����x2�^Ҭ��gf�q.��,5��W���`��n%�����������c�J��c�9�b˷C\anJ��=b�'n���d�l���ܖ;R�t�4c�A&�c�9r��jDZ�j����0g5�X��p6�Fk�0q��n>\c�-��'�=�#�]/�﯎�`/���u���n�ˈ�h�b���B��ݗ8�BQAy�u"�B�G˨G��k� ���?k�B�S�D�� �i�!ї拷�� �oՊ�#����K���eJ:�P;X�j����Y�,�ѕ�J���I�`��	K%Nd�7���W���wHo��^���i��j�K��K�B�����#�.vwX�k
f���M��8#<:l�{��4��	fK��q�0��V���/ť_}'�u���;��ِiV?�g�)|B!������F�z�h� �m�~�%���T�:���&AH$ٿ��8��O��Rҧ��$냻��hC��s��M\7����F V"v�N�Sg����U�܆���JeI}��]��z��(Z�l�� �m��U�����0Ɩ�tr7Խ�@F4�UmN鬴]�(ڥ����9�Ȕ��j��
A�$i��8U�9�K��;�7��\��Jf:�jʹ����|��lK*�U;:{�Ҫ_kr�I6Ut�����>~˴J�����;���n+9;��
v�_&but���N]�K��5��X���K��V8呂ǣ��R�w��r䩅CѰ���A�D��SY'�Ƥ�s�}��"�}D�y9�W֐�4��@B���jF�d@;Z������H�EPF�Ɉ�tGJOt�V{#�jxr1����qI�*��:!sa���Vn�AL���G�h�j�������&��iH�I��B�tVP	��c�{cߣ��$�~5@?<'��%�k���S�0�;P-p�H�6�3�o�0�4��)��i�
&�h�C\�p*��-���L2��2�l؀e#1�6d�:+,�T�`������ 2�W���@��6�~v�����w��Γ,�P��_�&:��jԨ�~Ð��R/�Ɯ�/k�K�3ke�oCf�<E}_��6G�ڨ��Ba���p	�:(��,%�TI��{��.E�D%���	�~��5�x�1���?	d��*eD[Nk���Ey����L�GN�O@�*�� �E3˾af�KRK�j�<�OT~�bl`&<.�W�2���s��30�XU[Y��B'���
�O)�q�Xw��)�[܅��>�X�З7�����<B��W^辟z\�U� �X-�:���E�ؾ�,dY��8���ĵ�� �*�y����ؔ�_�E'���y�ɛ<�42p�l�Uq�4H1Ĝ%XS@�׈rKd*~`<��i�C���5��I�t�ܛjp��u �����	�+8�J���򬶀d�[AN�&`��=5��_Y.ݎ[������� �:��).M=��w�l�ZM�߱�0�?�_]H"58�n3�a�dnb��{�D�asA\;g,R��P�w�=�I�L��>���r�-�~��oЯ�)f�A�Q@��&�2�kƚ��0w~I�q�n����Z��=Lb��.��VL�Q���F�~����jñ4-��)���XI�����	�E�7V�I_��B�t�3Lirc��@�d(2˰����\����1n�jmN$�޿A�]��z8$ (3:`�~9����IT*�.��t�������������5����@>�ׯ�L�͂%~�>b+��7C�&�K�7{���D�0W���p�?, ^������~��|�+y�U��(�D�敕�Z����-��s�z-s:�g��0Oq�?i^}5#D�Efh��>s�x�m����9����_kaK�=R�ԧC�,S�����
܄�t�Ѝh:Ǭ���\�g��6���m���{^r"���4�}�!���z�z���~�ݖ;�'��14s����PD�\�2`CX#~(�%߻��M=W�'F���F����}'<	����S�v��:�� �)A��r˖19g����% �V�>Pl+��3�A�0k��R����pL7����'�a*��ΖG Z-���߹�v�]vup�4� ���/�+,�\w���P�f�ޝH�QƒP���g�	�Iл)=����̖�뺔��]��pS�ec�[��4(�����\e�bg�z���'	��u��,�`"�᧤��1�J��.�9Scm�ʔ�֑�"
��Ks��h7�?���[ ����L�u�[���wy�S5$+�/e�E(:x	�$��0:���bn�xs���mo1(ן������.�+�h=�ɧ�b�uֶ�
�ʺ� �w����t��lAYyFJbj?�	-�:ܽc,hJ��˦�/��1C�y��h��y`������S�|����S����H���Y|i�v�|��^d�Z̚Q�点:��;��_��.�`Z���w��� D�Tv>*�~�N��+ی��KqTA��}2<��-�J!r���w!�"C����V�t[��K~�;�sĭ�X'9H^QJ��\��B�f���v��a���F��_j�*�����Wwօj�Eσ$J���ȃws`�'��H����=/�
�R�v����������
ަf����J����w	��Ґ2��"��ub�F����G��Vg�x0��'];ԡ�Ci�H'����W�җZ�o�o1��,�w�N�oG#<N�n�RW�������Nz_�x�p��2z�|+�1R�#��*)�6I�X6}-y���I~�顿
�m�C�h?9d1�N�"���V`K��*S�=}���Z�"V��!��[]�x�����A�ޭ��A�+;_v}���G?ND�