XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*rCs��n璤TP��C��쳌�rE��E��ޙ��ӧ4+`�
sj.b��Ga9I`�%c��u�x�I��N"�=�kt�نlP��_#�^O����&��P�[K���Z��~~�D�}c��VD�.��F\�
(P�\F=���^�P|f0�wM����ܱf�,l�r�Ҝ���k�� ���N��(��(�O�������e릳q��cOh��Z�M����r6��).uф�Ps��V⅓���5�%�hhS$,�+��M-�c5|�^���b���L�~VX��+�c2|��e���IW����%�Z���5��m����I�V�D�8K� ;b�����Z�o`���y^̡X���)f*��.	E<E%��� yV�4z��v�S#�yj���V��x9*v~�Mַ��� H`���qQQ��,�15��)[�b�Rwx��V� )"���O�ɶ�RO���(�|, Lf����8�>�J}�[6�m)�\.�I,�
�h�!4��̰�@O���99ƌ/�z�>(��'�
6:�e�W$�b���~�����`c���R�e�I*g��Y��rK!?����y�7��ִ
��t@1M����M�^������ت�G�T�v�9��[wo�k������5b�= $y�v8��1y�p�5�M�p^z��.Xj|���<ޞo1:�H{�0z3f	�zғ�Tٯ�h���Ԑٳ�ШE�_\[���[O�����$^�����d�dV[e�L}��?����XlxVHYEB    92ce    20e0�Q��0��\�X(���?�����b���?��~t�3lV_�{4!8/�|�j��z�g�����H4�4MN�,�j��:k?�sHj�Bݛ[����O˽���zh��y<2D�����Gg�~|Ր�����fʋ��V��t���[\?�V+��&؀>=n�bf���f<�o�s'I��v/�f/U���a��Wz�!�[���� 6Ϋ'��=o����y�(����ؼVTφg a����/6U�LԐ<�dY�T�.���F�r��4at-Q�2�o�9������4`�$��Bf�u7T1b��a+�I�����37,|��.MI��N��7��O-I7+�����!J0px헪�>hU�����p�nA�m����DWN��/��@��{���w�#Cb�l�ڷc�p.9Hy�NL$@���r���^Ĝ_9�J<N+���ɤq�v��5PqJ�XӴ\S&�OQK'hlO�L��8Q��,\��9B�������!�øv������1��]�H��x:���[o�:l����Vd.[S��M��u;��0y[o�{n��&˧�\x*�<4�0B�|7���֯�/�1�'+ڲ8����#����z��w��LQ�?eq������ 3.�cK�L�u���E�� �܁7�o��ԓ=;G�
��.���G�a���a�2�G�� @8��.\6<�w��+���&;�^R׏Qn߆	�QAZ[-7.<oOhc�->7,�E����[g�he��giG7��1�	�N����P:yR6Bn�1$I`P*v�����Zz O_�I)��s��;�2��b9Z-4V2AJ��v���������JtQ��,(�����{7��Jh�)CO����@���P=:&���B��F��4ms���B�}o�0�{`��3y��,�8)�&\����o�S'R�z�0)�kÒ�˜ !o�Q�'w1��Yw���_�B��ݏ���tݔO4EF�^��4��l.���@����b;za��/֋$�ǆ

���k��7�ᘏ���is��фw�݁��߿��?C'/㬦�u��XU8��؜m�ߜ��
��[�z�`-����1W��o�9q��
N�.�v����W������s� �?�'���	�!�_ce��C�itC��ʠj�%��筧c.f!d"��\��m6��=����V�p�S(s2HMWӓV�国�ZЯ� ��Ư�(����� |(y���u��NSDV��G'Kƕ��hdFf���sd��AW�ja�f�W�?ѐ!>�*��iu�_��Փʃ�N�Y��i�M�]�u�:��I�� �ͺ���{Ճ~�i��ٕH�-+�~1�Γ1_�є\w��O-�ꄚ�e��/_^|,�!j�]��8�K�j������o/����K�\!g '_:4! �}~�=�a]k�$5�A	�F��������%��X���7��=x��5�!��=1��s�^�����uq��̗c�ҜwO��S�Z� M�������>U���,tB:h��F�֒$#L��;�Oqfw{@wH	�2t(8�c�Y���c�{��H�l�p��]��l>F�w?�M�xq��zL���N^c�Y>͔drj�Jcm��=���&�:�JhE����!�(&��C�Nv^�;d���o�)D)�0ˋ����?�+߲�[��L��mT��T�dʀ;�r�9� �����Y���0�,����n�������q�#�T��R���1���BjӉ.O��+:��N�c�\9[}�����'C-m.3����Gڈ�7c�5R �׾��[���M[�эj�����ɓB
�JS����{l�+ވs��YE�ʚ鏌)!�~+����08��~>��E4?!�%��W�87�$"Z�7.�8��xX#q1=��&��kom�#Ǝ����l��r������&~I�^����J6jPW��BX���C�z��ܷ�QCj�0ή�V��Xk9�,�җa"�����1�(v��r̠�x��&Q��~��,ա�������ֿ67]�0{;�o��N���z�y �8'H?r>U�W(?T(������(����58r��)���tW�jw�7`)�-�t�L��P����9���4����%�fRB�},c	�	�����f�ٙ��,q���j�KK�p�IN���I����7iu 
�����	�;�.�T�#�MЎ�T���D���67�3���ۓb q�:!i�׈P����}b�ip����U�z{6�1bm���QC�h�02o����w;߮#�b�ZE_|M���A~�C�����S��zf'Ӧ�>�����4V���xr``�Ց�E�]k4���egP��o�����i�+@;�7k1��Q��|J	��>�r����1a�F��R�{ �ogG��	m3�O�| �k�߂��P�J���(?��C=��$k�`�Cp�M�_���j�+Ui2��z&+�[J��"OuP��煉Js�!��]�o7YZ��o�.}u1B$��+lr�AEPQ'D��A�-d�/��t�Q�#���͂��ݯ���/�vfW�%���2���dR;G�|��
�7�Z�a7
v��[���.^rG j1�Y$��xtO�ۄy���`��C��2B^����U'@ز�q�b�;M�t�\�t�W���ֲ\m��RFn�g��	�ȭ�1�Q����)�1?%��T'�a��t�s���#M,m�����y�[�.c�_����W��v.>�Y�[��'����b�׫b`�!�JI��f��:S�e�L�7nL�ˍ�ZJ���\q)Q���(��6�"�p�pft�hW]�:#�|�봊��dɩ]!�;�d�k��z�o�r�3�~�G���9r8`��>���]�Ц�V�2��B�],�Z%OO�۵0�H����"���*�&S�N��D�Q���3���&���]���m��S{�4�Ω�X�]>��*��o����#"�Q�Y��4$Ѵ|t)XҜ�_��Y�0�(B�Is����x�"ȕd���4tȄ�T60�w��*`~j M���n�.���:��;3Lě�dK�z�"�7PE�k|�0&�����7���4���D��.p�{7:��b�5w��W*Az(W
\mO�f������c�������KF��X��l�Ѭ!��(������Ƽ���8ĵ�Y��U>h��2���Vl���3���<M:���UA,V��J�[=jp�x6GQn �	З�k���'��2Ko+�]�.�6���S��V/;�>GU���dg=&�X_Pq́-���E��3��9I;�##IS�.WJ2��F�'pX7J�(������.R�"�ʙ�킏��4�(�l`�jT���	�˖Mp����Q��p۰��%��:��/F_�u	Of�Z��d���� �%7M���c�U��wdE�C�1@_�[�3��N+�o=�bB��b۝�d����H�8oZUf�%9��.�];�� ]sE�k��yF�"�� �jK+� @5M(�}��[2@o��g�s�@���K�Rgt�I��5��"���\˄��ӻ�i�����Q��h|ݥ��S��S�4o��F����v���ǸH]`e���.R�#����
��;XI�?z���]D�[gs�,�9�5����B��eQ�į��]Q,����&Stz��H�8�K-\o��Jj�#��A7�"HS�5��$�ڛ�Dt�`#�.h��Ġ� �E��Ja�Ss����$�&��*�V;�j����~�Y&�����HZo �n\��.!�f$K���}�d����k��)��Z����$�@f��{c��B�̨U��!�]Sÿ��$`ǣMK��޹�fc� }z���Z)%�pJ"�[�/��Ee�I�����?آO�Wy�W1$��$�R��e��f�#g����'�?�8vu��(L$���&m�Nl��F���Y�QQ�0-*of3*0�����c��MCb�#6��%�Y�g��O�Pr�?Ҡ�Kҍ�8ٞ��f��E��a|b;̺������9$	s8v��2��ύ�����4X��(���Ԋ
+P�1@s	^٨��W�7D��SlS�0��F�BV�-8���3Η���}*�:Cz�D����ܡv+�����e���E��{cF�%+H��ㆺ
�Mh(�ף��m��9&d���n8�9� ^VWm�o!)!��0���>���� $p��p1INV����4�'~ò��E�ގ G� Q|�/>8,��+�X��ī�(���������rl��yQ�A_Y���y;�U��b*۟d�1cH1/��
+��\��,j��J}���N�y�敓�#�q!⯲#�� �/r���c~��Qhk���N8��&�t:��8v�q�	?
{|D���l*.q �>��v�H�a��+&Jʘ@��Nb+�$�� 8���,�.��#~}�p��ϔ��#,�_<��fbR�f6s�1��pZ�|��I�¦;��Y���5��`l��������d����e�������Cp��eЇ�~2'�wm��v<N�p#9�C�}����틓�����	YpP���Q.5wp����&��GA�)O��s�g�ٌ��Y&��,�$᭸g4�vkHQ�%N�x�z��%o�QX�c�b�'S��y��v����t���̳�t<�#���+��W1��<�����xщeV����j�a������.;���Y>g�BV��������=E����Gw�W��S���:�r�J�3�]�d]EJ�+V:�Sk��,���q"��zD�����%�l��+0H�3*6�*Id��#�(0>;]8Ű����y�`!�a9�S��.h�t켴���f��WV�X�����t�Ce���@���wwrn,�=�t&�kJs���G��O�����bۑ��t�F[;\���,�n�f�J�-�m������is>��A� a�g˽�"�!�
NA{�O3s���/׾���%QEs���\/���:$���7�<5������������h���. �.�*hj[�+G���nn���Y�#��l�@�P�}Y��+R8��}ܸ3`�����r�p	)6ešu��`07,�]�N��z��D�wXF�w��x���	"h�F3e�K�H���֪a.�ͨ1�w,ӂ	���Ka���t��Q�in������uj��$5��!<N!�h?%�S�R�8(�cU��<8�˷�5W��&�0��Z}���`�~o8.A��LOގ�G6�@p�	�3<��uun���h�L(��9�Y��؍����'�Ayn%?,$f#΄9r,��xxٮL����@Oq#t�>�M�(�􆃑0�|0ʓ��$��D5 ׃��q��Ť�3���3�M�g�]x�f�˾�ȓu�$����vcՙN���m��=� d�%/cIeㄞz3Zʳ�˥'�\��HN	���od|,��*����}�֪t����[x��+�f�S@M�W<�u�`�<G�<.n��x�Ѱ7��Y:��l��V�&{;*n�G�jUT����s,=D3;Ur~�@����*'<�`���b��)�&�s�0��&f�0w��Q�6�#�2����|�₪�hI,O���XcOS�7]崡�;O�@�p���6'�p�nɍ%*]6��2�*�$SU\�J��s*�{S5�<7]9"<_כ�!��g9�s����a-�͡7����c��w�E(#���W.ol�^�+f���x���<��!;O.��x�ҵ�[	HӇ�ٿd��+2XP�Qs ����(&ō��ˀ^��}XC�{-Ŧ�]Q�����t�k�\!(a*�?��N����u|�U�������cG�s�j�S���s`���z����A7c��4�h��l^Gkz���^���.!?�~ɰ�5���ר>�.-tq�Gϋ	�Wn��c����øc('���6(f^mN��T�ص��5�ʲ�g����॔4�9�QB�|��z��L��];O9XFR�y�6�\Y�T��ƭ#�n������v�zc.�-ċ�#�lA �}��>�|ɕ�Q�?y��~�X���Y����ay99��sC���ϩC��x[	��"�I�8��|Z2���`ww�k/}O�W��Z��IL�M8�.�*ط��_b�U`�C/��I�P\	KWM���߯�F{B�;�S9
Tޑ�lglѼ�s>�c����3���*�Y
��u�b�Z
.�bi �3'��0����7&ttP���J=����!Kv��� d��
�M�`�@�L�Aa��Cw:�6'�+�srV�����K��hy���ƈX�!�7.X��@<��*�\h������Vv�g+���{�`��Y��p61���g�qḩ$:�3���AP킐���!��%����DA��Ң��5&w��OO�a���,y�m܎J%YĂo���+A}:}�ϱ��(�b�H޶��֣O��f�n�6�*@��MzJ��*�<p]���߱'7G�� ��M!Q�X��v���*��&uJ~An�Q��"�B�p�JZ���H	���S���&�����Hݠ�1& �S����ԼU�2��V��h-��C��T��#gg����M{L�yr$P�A��"+x
M�m��~��W�T���ﱘ}�ܝ;E��F�p��"�nھ6a軂�Xsks]�c[�T��ñUz��/T�1��Ib�4|��R.0,�?Qc��3%�hx%+�V�}�r)�*A47�~<���k÷J<���0��!b��aJo�B	��~�4ˏ���d3�T�d�%")f��w=�H�᣺B�7�j��Ǖ$�ƫ<�D,�1�H�^YV2�"����X� I}V�*�����3�+h�*�V�GrO����D����k��#ae�&� �ˮ�m#���h��N|��ljf;�ܡR|@Cc��N@>����1��క{����A�8��R�1�9�A%:V�;ѫ��Ͻ2��.nUR�:y���a��骉��Z˘��nX�y*��w*����cH�_	��(YUe�mi�1�C�@��y2�H�9��������%�Q7L�$@�	��^7�l��<�5]?�&{դ�� ����A�1Gܝ�l��%4�����*�����F/�ea�h�$�j��	�	�F��< 	r�E��&�:����~�.(͝�S�`?:hQ�������y,��¾���/��1fZ�en����n(T-���2g-]�O��`F��h�D`4)"mrة��/���'���;p;3=,�f��?���R#Y���\���#'�s׮ұ~V�\�]T�0���Oj�1]r�i�6�L�S�g�5ʱ���|��ΐ�p�c)��g�An��c�w��v]�Ϟ��Jv`�v����mtӞ��z~�D!+&�V�#L�63�SD���z����y�=҈c'��g��q)5��~�@�s��q����D��?�R�)����s[)�De�����guRWV���Dd)M}�ڍ>�śB�ְ�Bf&c�R�d��<��s����ά���Ai�7���yS�I�c���c�Ds�8ÙXk?	�x���)��c#�&m��+lP)�v�R|a�J������pk�����W6d����E���l�M�������5�  ��������mE����OY_F��F]������c͸ %-�L�]yy_����	��^?��fd�!a�v߀Gɝ- (.�u�H}�p�f��LN	�8���'&L���u���7�Jp��m�u<���M�Z�[m�� .��bԪ@�	�=��?:��/d�<�� r[%�xf�֞�t'���Z��' �o��[L\v�c�8ؐx�H`!9q�������"=�,��^�[k��u<Z��F�7����s���nH�o�0�`��r#sy�:��Ww�檢���f�U��y�?[b��E��A괣���!?��X���[�_�|6�/��up�x�t��,n
e��V�5���y+w#D��R
���{�$��6r�FWML�d��g����:H;zv��f`��������043h�J���W�Q@�D����;���s^("�/�B��@���d��꤅�y]�x�M����hZ�h>�N]�*ο`�x��W� ��=i8%��u�mJ����͖B�^!�XN儞G̃l�>y:�c�9h��ف|�$����B�m�Hdx��C�$q���K	5�Q�9�LnW�:Ԕ,_�һB���ٽ�X#�
�ЕJ)!�z�9.�/��n|@�06U'