XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Mj�Ҙq��5���+��I����@b?dB�v�����և��*��N�̐l��c��VP�d$v	=��>�*l9��� p��+�$����s��t�!�'�uMݞm���S*)wP��_)���#C8t���=Z�Si+8A��l�7ѧ�~ػ��V^M���&-NCdO�H3��7��f��Yz�qH{�OG�n¶�Sr,J�]z7W�06%Ak��nI:8S���i�Yp��K�y$S&F�`�b����E=�gV����]o�m�Kņ��y��hv*��[\����u�[��֗4Zy"j��_\�C\��<�/���.�yu!�d���l1��*����pY�E] �m	Qo��0�Ϩ=@�li�׿�N�$ϰ^�O{�&x��`B�yg2���v����;}�٪߃�o�$�����W7��Ԗ�\�x�V���^��m�>bj������sk��&׌o"�+�s���{)?�r�)��k
"־V�n<�t]N7���,cF儠ٻo��D��c���'���$5���B.frp�8���5��8�B/���U�p��ODѹ�@�	�V���W��>|�Պ+��&�����s:�	������IpJ����v|iPM������d�[}ʢ���*ֈ���ona�EV}ڜ���O2��R�ϳ�߅�F.ՙM�b��r͛�	G�Z=�����&
���K���@��{�k���y�Ĉ���"T� �2�bZoqt���������N����-�_�Rn�|Ԝ[�*B~XlxVHYEB    c227    1f50�
�K�Ņ	�4����I�@MI�"���*��so�%�̞�Mk� ��:�? �4����;OZ|b6aH�'%1D[k���-��-��w���D�`���ɺz���{r)��P``�IR^3�������@�[����[���m3��;��0�"G���X�vڞi�g+�[V��96�c1��+�=�*T���aAϼ�ߓ�
��A�k����aYo��*�,�̚����P�k�֊ү���.���Τ�� ;���H�7��P�F��+_��f?OMZ%�듋\w��P�zt��{1�T���E�¡R\p-!�X@�j>:�����e5[��6U�_g�@@���� �JC����,��m�M�/Tj�{DiT\�Rw~�B7v��T'�MR��BJIǂ-z����ۍu��/� �R�*�!��b<hX;㏠�������Z%s��m�׈�TX��u*���C�ԫ�2�߿M�� ���1p��ӗ�!;�e3\��@��1�P/��0ҕ�D�k5�@��<v���2�h�����J3Ϋ=�6��3�jhY����e��UP��kJc&��v����K4B!�T2m�ֽ�7KQ�w �d3�w7H
"�+�v!��C��t�ơ7��=��<��^�.���"D�m�����J���ik�x�\�M�T�#��`��� P:ޛ# ��P�ʇ���+�-G��#�����>��޳�|+�ޛ� '	ב�1� ���.�K�y;r&ꊤ/~��k���2��f��N�wOS�����%>�\!X�\�]���OX�x���NM�~Cj�'[�Vp�법��z���f{�B,�Es��u�]pJ�f�W���*t�B]b��C�ט�¸��͗����
��1�'~���@ID�IA �F_]qz3�0��=Z�����t�/�O�:�1��/���h}&TmR|_�w9� ObPߣ��sG�7�HKD�G���^�2� ܠj3~�ٍa�[E-ʫ眶`x�G��0��M�o��H�O�����,� ��������՝����^����l�D*��j���������_X���O�RRw��%��I�)w	��x^��E�T}��P��i��GE����JTx�Wݥ�Sr����i"�_�k���TH��zs�v��~�}�}M3/f���QϞ���Q ��QS���z%��O��b�05�TP�G�w�F�]@�H�iu\̷�!}��S\��G.^��ԇC��K��O������v7�G��
�_�R��I<3���\$�ө���� ���K�O�)wѺIj�������c��{/�пG��Y�.�Tׁ"+��Vc�����iܪ���3��e�L�m"�e뫆Z<�eÏ/D��Zk���y7�@>��1"���M��9A[a#�����&�C���~g�>�U)�UQ�Xu��+��5u��s���ݡfVʅ��RD�`���u�2�l��JR��$���N����J_�HpY��h�"y��2���|�0� n�P���5����_��q����ǂ/ll-M�A	�C�8X&M���$�(E�������cd�K)Drj��ϗ��x��ސC� �I@^9#m��XU!$.��!���^g��lZ�M�%o�VK��-sV���~�J~m��0?�[�m�{���W�&��>a�Y%J��mp���(G�t�K�*|�0�O"r�d�C-���X��3�i�o�A0�H���
��]�Lh���$d�.�����ګ�g��8'�����f5� ]1�|.��>〷�pS����侬^߼��(�W5�焪Ժ}q�2�ӵ�L˝w��ǻc���ܥ��:4!	eJ]�п�1��-�O����]�m/�O����Su%�J�] ��������FC�k���Xc
��0۲���{TXB�?;G�e�+�}�t85�EC�57�
o��B$
���
6?��u	�g�� yr��Ϳ���oo�$4��R_Zv���K���.�E���*-�|��ܦ/ˣ���7����݂/�H�z!0�o��G"X����Km��\�@��8�ͮ��P�~e
@�=��U@e^,p�kz�g�)���䰬��:��b�UA/�)fe�K�
�^G�Ǯ�h�=�����#����dD���R��2g���Ƶ��ֲa�Ш������3����>Æ��kY@W�%�g��n��z�������p���"�� z�N$
�j2�pIQ�a���}�xF��`&����\
dL��ew��!��e�Z�L(5�f�p����������c��+[�Q�+�݅u���yM�ܽ�w�Fsb��n�-Ko��9���^��IO+���%mb�F9h�Ia[�X���,�>J��;>�\Nv��P�l�&����1k�k!($��Ȋ��]�**�%�Z7������8�����H5����*����:V�ǂ����>0�&�E���y��5v���k)G;��)D��K��"���]exm_����X��C��o� ��%{�mMʬu�%@RY�l�^3:(�J�ʽ ۴i$=�\a��	�&kv�|!�~x��8|��I_H�J�Xq�"�J~�k,�O	p�F��k;ԡp[�>P��g�J��N{X�i����l����!e0c �@�MQ�[~e6�'8ޘ|Ű���w����cb�m���eԔ,�]��$���6��Iӫk��R,}$�m琄��\5�Рw���r'a���>��;��]֊���L�\���%a�.A��oDH5�����'�\�-�&&Ԑ4�+$���f��i��/��"AЌ�H��rY��	*��QD���YD�kR�_y%x߳�ºd��T�eF5�$�:JQ��4j���F��aCM�nx�<����	^�����g��.{��҉e�f:&]��L�>�R��"�Y�b��ο!�00�Ӏ�����k2��3��K��_85BĢ�,5sO�E��|
�h�����������E�{�R)qx`C ��q���i���CQ#"��Sg�]��m{Β���6j���]� ;�	�2�?��q��#SU�td�"��;%~s.�H
,���e)�����kg\���܂@W��#�q!�V18���&���!�@,�ԨM���D���q���]�9�l��1O^���лYՠ�x��G�^o�W-���Z[�3���QR$���}q��}4��r�-,�#c-z�B}H��*~�.|?�{��8���h~��Fj���y��+D��֑39���g�?��	8c�Ψ�����a���;5׹��T7�r�*�0�ڼ_Wl���8�U�B���%*f[���3�t�n�1���ѽF���ħtvw��((c�.�q���]�C��ҫ���R,0�|����.��3�x�]OE9-�2[�}$9G�R�*I�{;'�<�����L;�u��L'�h�'��ht��ua�mg����
�3_bUf�$Ia�T�l������_��|pS�����ɒ�7�R����r�As��^c ��~m/_-f&�֓�u�7����wN���@�Lrbl�W�?N��w�F�vS�(��#[q_�^uGG?�ϕ�~�W�\$�����bw�ݾ�����8�hy��ٚY�v�(����}W��}�?>A�������O�7O&�Ǫ�W�ro��pH֫$����-dF�7�P��\���ܧf+�O	~nw#����;�d��t�x��gV�/���K��S�
.����߻1�>���;V���vd�)���RMu��6\����0���Rmy���sa7IE+��}?߬��Q�ѵ�� ���7ʿ��H�;x�~����i��{�(:�!�N�KP8��O�9�I�u>�J��lӓ
Ǎ�P�BB�*����ʝ�Uj��G��[E-e���<$C�7<��^�<0�S3J��F���T��-��M��o��Ua�pL�]
��<䟊Gx�����e��=�%��b�޴/��Z�:��8�㵃��EB;J��JN_�YrެR�:����3L�Wq��?��&��|�a,&�?�^۝�8�Ť=�2�#��R>�յ��/����y#����C�=0O_ɨ$u��2�^_�$O���9N���ċ	��wu��W��w(�fm��^�C�>���(u��P\�`�Ɖͼ��O9H�|��k �FOٔ@�(W��U������9�e�K>������<3�0|a��^�h�DFaY�Si��z~^[,H=�������!�K-���f& ��B>�{���7� ,`?v���d�JE��Դ��h��%�t�ڮSeM6+tfѽ2Gx�4�H7�p.}�&֓�KϡGڬJ�|������U��0���O�^�]��R783`��Wa+q`-ȉ["��5��'H&)�b�'w�))~�:�Y�|M�ޡhi���7v \����r�����AQQ4%�1����]��:��Jݦ��JQ���,����B\"{�uY�Q��y���ȘQtU:��b֞�����([�_�u�i%�7�l�%� RT�e���Jc�M�ex�'8U��߀c�Q1�30=4?�eI˗�h�0G^�qi)\~�����G<���'`N<DǰD�O�Ce{&��XmD�z[�y$��b��$
,��w3�ʻ���T��}=�6c4��Ij��ryk�m)����m�ĝn��Ҿs�J*���������#��@�������ݸ|����f��A��^��ُ[M��%��L�7��grȰ�"<bI����X�����O�*y���v���`���%�Q��׃�ư��)�s�^Â]����r|^tғ��\R�OX�?q[�_����%%J83�H؍�*ŏ~��l����qg�d��"P�'�7�Xz3�:e��,�^0�c)�T���Q��.���}����F�*�M�5�Jf�1��na���ydwq+��tA���S5`l��z�B>�ճ-����c��#��1H�=<�R��J��-��A�1����{(�6�g�r
��A���@�P���_�f�`�7o���f?�^��=N�G��H�b䫛�����ȘIN�ƭ����1Y�s�}ǨP+��{�����KvE]_֓�bf�dm/yĥ�h�1�rQb�Ӭ9����-��X�A-�:�A�7ͧ>㝅ۖ�`�\�2'��I��8�g#�O0�ej��̧����]}��ї�HA��XE�3`�VY�ΐX���;�6�"� ��f��[L)"h��[����5S���,�!�?M���zMjj��z*cfayz&��Q�*��ΐ�%(�}��L㬍���a�ٖ�j���to<�:�y�S�ѵ��83�ynS �����-�*�:�KTA��ǜ�-�͵Ķ�5O^i�`+_R��jmp ���6/h����)x��C)�m�!�h��9�̻1�9ǎ
�su%��+S���X%ѱ�q�j9P��C�M�qh���3E��$����+��PR-��LX?3|�s�h�t���^�mt�����r$�����4KPg����F��0�҂���a����f/_���,�'z�7�q���9��H��������Pkw�\m삛�[Z/��zT��+�b��
��kd��P�P���[�C3��|!;��*�Yץ�D��9%���иM"J2Q����D�"��%։W �p�����w[5Xp�kκ:f��b^���g|�^|�H0��	�귲��c��h:>}\�˙8�o��YB�˜2�DĮ��=&������OF���G�3���i��46�#��لp�r�>�\��9j3�7��n�L� ������b�>�Y����W���7��K?�cPz��Կ�XU/��VA��'���v4�����!Н��<���Ͱ���,zy©pGwV�B��}���E箵П���y����!z�-T���D�����V�s�)(��E���4�D�*��_i5qBdݰ�����F�\.��?����{4,'��J�zZL�C'��ڔ�5���k޼��W�EQ�
���cE��?��rU��;�����5�#�.���X�lħz�rc����[����^�^�Y�C��+�0�Je��0�/�V 1��W�j���������Y��e<����>��C�r���k�a�_r�H-�o��0="��4�=xت���/&@��X6��} _«=�,h���=r�B�ާͅ����04{�{^����zD�dG��b�:�.�!�~�Rq�h����GQY�|�Vjp�ԋ��h�q�{Z��$��gB���n38$&�$��a.�i2RX�q�)s��M�`�Q�� ҕ�(�D�G$��-'������<1|�5�ޭM+�3����<�rF&Ns�&q��z~��&T�i�V�58ƹ%�>!���}��ۥhB���Bp�$oovS`J��y���]���� �1+��9�,*E��� ڸ��/��GN��NW\@SX��8��̛��#�Z�o��,W}���/�H�����p�)D��#�[I�$B��heJ���M]w:fm9�`�,Ǡ��1�bBSq�6ڬ?c��5d_9�&l�j��8�f�B��A�+�?�P8U��d�{5FHx�F8�#z���-�J�D��sH���I{�Ţt^�:����w@��IꈅnE�����j
��%����tD:tfr���	fʺw\�ʿ5�+��
��Ud���ʹ"���*s��(K�3�k��K���^������p�N�)���J�՗�O,�Z����Gz4�xOiꋣ�(�ne���o��yH�L��䤝�f�i
��r��<����w�O^2s��l�UҊ�w* �ނ!�M0�HH���F (D�21m2NFP.�7����_ �:z>���������aq��Z�0LmF�N��
�K7��#�I�`J�F���2��i��,���� U�03!�S���*�}�;��Q�%!�hO��A븦�GD���kU��]J[fp�>����K푛>b��	�a�F9���j�"68n�*O���BA|��@��?�+r��}�u?= ��}���a��2~��П��5����K�^G�6] �5���
R��
�Vr=B0=��ܩEg��Ԥ�����$sF����q�`��pp��DN�mKƫi���@"�r;ЕĻ����<��� ���Z|M��[�x|sQ@�aH�#iLG��87d���f��F��b<��[n�mܖ�"����w���i^�����	#Ǧ��%���Aգ�<�R�|8��/����E�јp�{�·�ł�۝Α�B1?�7��R�Pv����.nu,�]�~�����Y�gP߿�*�e�dL�t5�V�z1ě�0���O�=�eR��'�\e�<$c�޷5�Y�ڽKE"A-`���ի;��9�e��=
�&�!�WF1���Ϲ
=];m� �7ڋA%ԁU�A`EQ��&.I�YK�z��n.�U8�鉪陋)�U!��eBT!xo���(�zs�oZj�2�]KN~	���X��K9�R�������a��ޜ���P�)\��>W����D�����B����|26p�m�˅�ɕLE�~y�ٟ�Մ�l 1�)]�L^�Ue�D]�#	�u�,�G�69�Z�E�}�p����������m.��w�?��
Anvl���#ǫ�eI�#���A�t4秮�K�tQ�Ԝ����-A%3̕���ad�k���
Q�B���p$Sj.e6�)q��p��CNnU��a���=A��-D�`�90p�p��dB���_������=1)L�Q�ۂq�8��������	�9BB�MTxT+��/�f�뉶6���)^ 5������+#��5�$9bO��O��=�݃ދNu�L$�cK