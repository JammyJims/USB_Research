XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|�������ɫ�G��d�C��V��V���!��_/dce;�r�0=3<�z
��q���D�p�g�1!���M��Dx�F�;EY�=m�M���=��x3�8����^Ӓ�1L��0~*�����V��s�1o����C�{����4\A���92Ԣk��iK{�~�;¯�@D¦�Xh�v�sD�,dO�����<�e�����-HLx�̖'a��:�����BL;(��Ɠy
o�\h���]Ԭ���-��
7%O{1�����٢)#�j���x��$,&ud+Y<L"��0V�`~�8/�/þX�R�^Č�:��q��Bn�ƻ������]�[_P3���g�j8��ϸ�i�m13���������`� z��n��9T:��'�^,���12+�����'Υ�p)zGƄ��u�r�B���D�ۯA�KW �d��+<�es�v=�R��_�1���u���7�_�R���	Y�ì.�����`�[�������0��ӯ-�2x�I7�Ciǟ��
����EI.��B~b�F�P�ݡ3N�s	p>(���^-l���!�@�A����g�1/2%����z�cd���	��P�Ol\�PS.�dE��V�
��sz<:���l��P4�9Q�pF��)� ��v�"�x2>QXh�~�R*��|��F��Xx+=8��ͦ��s�ws>.�sճ-�۲�f�2 2�ػ���)OT�ߩ������69�	���u��Q�;ٮ�nD�Ǻ��=�XlxVHYEB    6dd8     e90z��#��MR��r?��Xb&\=���8|��1�]�h�d���Y�+?�1���4�eM��]�'Eb`l�ٙ7���s��z��#_b��֣>��9s�G.G#JT�Cye��E��7:�3�����W��6k�+h�
Q�ѷ�����c|�X�R�(y6X���f�~n���C"���z<�ͩ�y��&l2ҍo��1;���*ԍ�/��~*��R��hX0�2_�Y��>nے�LT]���e�F��|��E#�`,�^|��^Fy������O魨�u���l�yh�`�=J����D�e�0�̾t�v�A�����O�\��5��U� ������SK�Qo�ŏEʨ�hk�]��(?���V�+���׎�/^x
�����,�!��%M�_�qcA�4)U��%0<X�?����«�����Q�d��s�loR{��)�sT�<�QI�����(�d�qS�վ��q�sO8-��^���w�pV��T�H�5������X[�Y�8W���#�WpՅ���i".��[�{�Y\}��`��}���^���b���B1������C��v̀��zz#;�C�����k�se�-q�2�k
��a��i��&�Ū��G��}�G�o����ij�e�O�����cF,�2���y� 93���v���ѷ+Z�Z5�4��^g�����K$Qc<�Эi�⯸�wT +�޵'@��������v�`�$�`V
���s�X;�05s�~�KlX�	���h�#Ӗ��&��|f��O�@�����1�m������܊A?"�*�p��z���d��R���^�8 S���K�����Q��=��s�© ��bwP�i�i-�{I�w�T�W�8�K����� aa�N0�ty��<Q1���x�Ι,���5eu.L���*���U[��B�ά���J�s�&u��z�l-�`9C �-kV�GY���B�M�K?e���:n�I��wl�-D�^�l<8j6��'�e����υ\7�rbTj�RX��'���00�וt�e}�XEE��Դ����_Ǳg�v.�G�D��xW�6�Z�t_���j��i���oMTj�C��(�>��P�ϐb_)��U3�S�*N(�;XfUP6�H�'XUZ
=�]����Y���,����&���'���T�dM�p��5���edcU��P6��Tڨ����o�������GjL_�ׅ?�(3E���Ϗ��k���y���3�abX7��V>m�sB0�UbAf'Ǎ���ǻ�1�R���j��m��-�">��:.Q�)���,�m�f���<��Ľ�F�T�2j<N�z�p�[@�
4�Bg���zb���V�R�ҁ1���<�����vhU 6�����s����
��m!)^������&�o�]Tb�})E��S��f� �����Kb��,#l�2��|��q���L�u5b�X�*�`�1���g�f0��J锿QHƢ��?��l6�r�G������]cR{�c6 �x�Џ�
��؏i�3�cդ�W@�6hz=��
��
�k���J�d�4�毲!��8����O���f�p��@ǹ*p�%����R3fYjlpk����ad20���$&m"qy�h����J4
?�3��0�2�hme��Q"=5*;� �n��P�D����O�)���x�z�,-�)!O�v+��
��p�g�t��O"LCp8�����jQ�-J�E�x"k�/���2Xn�o�
_C�8�=�.w�\S�5���M*�Pi��.�˘N�2�����0��IJ%�fÄ䅠�.�1_�+k@�)�_(��o$秖�]�Ye�1"ŋ#�ǩli 47ʂ�9�Γ^)�=��w0��|@q����AUY�������*����4�����1�n��㭹@N����U�*c�����%�B=f֯<���PI��$@�HfB#E����-���(i�|4���봚����rw���F#s(k�Z��m�vb5��&�K�-oSs���ЖJY�)�%/Br˿����p&�������3� 23�7�:
�T:�����w�1����[���tp�(����"���vu��8���ͫ�c�M��-����&����sد'��J?�O��v+�Rh>�I�����ͧM?2�q�me�����x�v��6$��f�FG_ј$����׿�G�C~Z.z�5u_@�+Ϫ�A�'8��Є��y����ͱ��|�@*�9*�d�0����y��?;�Ñ�(�X�J��R��kQ �&� ��V1d-��z��ّp����x�X���lG�(��#P��SlFw~|�Ǻ�Bh�h�"��Ȇ�&E��_ hQ�w�_ �2�'�1	*��� �}$�2ё�c���F�A�e(�=@'%�H$>��Ϙ�ZqEB��g��o�H�[�ͩ����9�ԏ�oM~��oY���K�����t�*�=�kfd�7�0ЋM�,ee�	�Ϧ�;�٥���T+���E�=��w�6ŒT,�s���,π8}���7��7�nɈ����Ȣ%vj|�m"�f�P26�a�:3P8F)�t6b�tgњP�������V;���|��@y�{A¸��^�զ��I�P����Iwi���u��9\������������%�r�����KA�B3.����FcG��W��-�BZJvj���9�C�'�0�w1��_5�B�X����0*�L�іtR��J)b6��ꉇ���9���NB����>�d J��ۮ�Q��$�_9������7���BЂ�g�p?�*.�T���Di칱��]6	�?�G��P�>��#�X\���掰y(��N�c����?:	�v��S&�'C��K��q��\�˅#����w���qh�K�m_1*/?j,ڂv��o��\@�Ssʌx
}A�����}*0&LJ5==|���:� B`�H%r�/m�'��s-L�u�7\�#j��9�y���p�=���Eѱ���A�H���;/�Q�,��C
�Rb�#�C��Qi�U�3�=�`6��J����c�!%Mq�^��1��x���g`�?��;ai�t����Ա~���9�e�cp�U4B�y~e+��# /H��dK�T~�E�=��9z_�Q`�Y�6��J/y�Ŀ'Y���qF��dg�VI��4C�K��{�;�Iγ��\�O��R#�/�]�M~����"�2���E-`��/�˳<{���s��� �Q��&E�5B[��'9�N�/�ۊ#���Q��p��Mp�4�sQN���8��k(���,Qe�*S�OF=n�~kU�:D4Z�(8:�֠��"W�}<���.����!�:�M�Р-��u��Z�r~������$
r��	�B��ªu��e�˚j��F����U���*w�.��R-I%�lt�4�~�t��(4=��<��&��Gޟ�+ϥ���YPг3g��w�~ӚD�f-f�EY�-xĪ����g���N�����4_���̩�a�)g��HB��Zjr8S[Ы!�O��Ə�bR��P-�wM��a\q����D���VUӅd�4�S���VG�9���U�n�I��[\�s˖�{u����4?Hc�@zU��_
�߀���lq���n������Gu����џ�G��e����(Jg�j�[� ��`��Qոp�Oc,���d��