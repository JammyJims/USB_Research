XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������t	�T�n#�
��r�2�Po,dt�E��ȼ���`DPf����w�^"���,�1�C�Z{�R���
���9��� 4���Q�1&��U#�C�&:�6�DWƾ�(�3X���ѡ�A?�=�c.��¾���Iz4Z�S�@V��j\�m� a�c�t{o	���xbq�pg��t���O��Y2����Ǆwq�5�ݭ�A��Q����稣����/�g��yv�^Uw�E0�߽Yڀw�������l�N��R$<�����cmF�j�����^��Ae瀨v��2Q��s������Z(G��0 @���ڼh/��Mm7W�\o�vrX�f#."1PU�>�}ľ������ۭMṣk$3��w��T#�����(k�����=�@F�KD���u�U�2s�B�.P6@2:Z������"%�%5�c�+��	�t�?��K�5�g�����Oq�2��W�ģ��AV�V`����/���2�W��H�"$G�����AU�	�t�c���vܼj�]}H����������@>�G�3�^ODǬhgd��{�M��z}'攽3��Ite���	���Ԗ��B������RR��1H�ׅ�m��p�Q��D���-�Yg��(������8��ƹ��aN,��#�UV0��_T�>
���-���H僿�0�*�m'���v�������|.�����[p�?�?�(M��x"��P �b���k1�Ӿ�npT;�㞙:{��XlxVHYEB    2907     cf0/��~Lh�f@m>1����u��.afot������
x�K���o����H�R�t�0j�i{E��?���x��5��eS��i�ؖ�Q�U�`��XG�I%Q�T�������%���W�/?� "�ɸ��ǳ�Ot"�;�U�a�͡��RR�Zź�W�Y>m0s��/rä54\Mqr����T	� S���zD]|�j� ���+�M�J��8*�&���GD��~�u��n�mI��:�y6|T�����J�5�W@��Ѩ�����$�_R���@���:�=w2Q0&P�L�Ե(����
����˔�.�݈��"^e��J%�4&�W�mv�ҹ���2�"q�؄�x�p�d�Z�9l�=�C]���_ 5�Ǩ�o�K�������_�j�i�M��DG�v�Tg����CBR��p�}���x�����p��D\?|�P13�%��N(Y��h��[�;q�΋� �ww���zt�$a a�U�#´O�gҶ�"�C�� nИ�`������r ��֓<+���R%b��Aa&�mN*��i�E00�}yr<��+}R&ؤ�A4{:X��
z���e��?��m���Hv�G	�[��?�R8w�3e��<f,N]���LH,��t����q�Gۀ�uF1K�����U� ?��N�+5Fk�^9a3l6�:�C}���id�V$���c8uд�Xc'���3�Ge����r��7?+�<���k9~���t�X�ڛ1\��,�N�Tk�+��T2\]������&j�C,�AV�v��t$G�h���<j����l��%D��X��?Ϲ��[��P5����� �gf����[k�ƍ���q�ޱ�?:�o7��t����<t���2�~}����s�����}`�<�ϼ�|}m�OC��,3�^��R�l��n�У��_=p��H�e1���_:n�}p7�L����}�P���
Fcj�O�RP6�K��%�� '� f����Ċ%�4�
f�@�!|�t�bc�<x=��2�2bA�I�H�A�SA��ǖ����m����[L��Ҿ�.�җZ��-���R ����ko��<J6�ʸV%�Д_�G�D��Z�4��U����3���j�:j�w�A���U �W9*�%Y	- ����+Q�ot��@tL9B�ٷ��L��{�}�j���[���uQ��y3�4��!�Q���b�t?d-��n}���s�����&hP�r����bg}�V�!ܚ�a)����K�k}v�n=r�t�{�˯�B{�cf��<��i>(F�v�8e�z�,��A١8R����P�ܙC�9�r&`�A�	C��ғ۶��9�X/�_@x��h@���2 
��9Y�n��])2�G�����}� >��AC|��xV����b�� ��j���'֪�K�zæ�1 E�H�ĺ�8��pG������s�{"��+�~�x4�� ���/��)���q�1Bg����7��PP~�T�e�[g�ݸ-S��8^�K%ީ�G�w/�l�eѕz�(
L��уz���9�U��5��3s�\�gk W�� .�uRm���р"�r��d�r�
���/�����S���x�ť�#[u#-7�2,+�?��N���	-��ҍ��e��Kc�.%�3ie$�E�9^c u�8a��׌�8���+�u_[�\�i��y>����Jhj�H®^u<�	#
g����_Ԏ���~ ��������܍�Q���vR|S�`3�#���g!&��J���=�~BK�Esςw�(L�A	�h;F��JQAj~pP���.����2s.�Ki�窉D��՝�����xj�!�ǆjd�1�U� `���tm���ˈӝ�F��.'�����x�O���9N���"��%����B;MfXrpVf7���OJ�|T�Q��ysG�wi�9-~��y�ȅQX���4W����*�S�����*���w�Q�_TBG��%�d���tS���Á��1�\������W-i��a#il�ВD�!�Kt-xfǅ�	����=zk ��^�>p"U[�`���q�8Stv��(��M\@7�
��R���tM�������hl�+M�)L���#񘈼J�R���kn@<�9_�� c6�%ǋIJ:J~����V �xl�h�HW,ߜ9�����v���}�܃��m\�#�!>��z������.v�x
O����2F�To#3T����^Li�0�a�$���5l�Q'O;�-�8�gCW�L2W�W���_��M��en6�����\�����)�������PڭU��ػf�؜�S�~aS�p�3m������m����$���x}	�:Ɖ��H���:k�����Ǥ[	s6��ڳc�#�s"U����c��t��x���F%s}�f��R-oM�]����(�l��Ρ��\a˗Nk/���Iތʜ�>C��_3�C4`��%0݋w4��u��[�����3B����I=�J���v���{i���BwUs>.�~0N1�����"����{A����j���4ֱ�ջ��\d�N��ȷ�Ng��F/����eW�nN��2�/�N��&0Gpۓ�X�<��%���",v�?`��$�%J)R�H�u���*�?�CV��g���]e��:c%l�2�CL�q��m� A������*��M��,��G�(X�@8s�PnW��g�$��W���$T��;��!�mx�p�EjoWyg7n�@l�J���y�(}#sČT\�>)]$����I���b��P� ��Nb�\��%y����C;�ٹCڄ�#�L��Y7��T�L;H��C�˚���8�>��]�����%Ȭ;��}hq����<w��J+M̄��{���:{H�dˤ��r������L@+a��?�@%��1��B1Zx�S�ϗ?oY�XO)ˬ�K?���Ha� sSFu��l�.��X:~��vK���s964p���(�m�E��#3�3�q���kuI���MĄ� �g9�
ل_RBMNP���)ǐ2�,܁}(�k֓z��F*�i~f���Q2��O9a�xO��\tT���:�3.�5�sȘ�2����E����&Ώ���~چD�B�'�83j�U$��B3<$)Ŕ$�kw�L>�7�,��zR7Y�) �B�.v����W���' �Xcup҂�!%��Ǧ�z��o�Vh�d.�\A/z����Gnn:͜��X
��b�fU��.�Nm	���06