XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@� �/up�����߼�k�=$^��P�`���r���Z�N�����9T32�H��6ۚʈ���[:����~�	�t�X���Ϊ!�����@kF��I�Ż�âh�1kzw֌R�Ip�.\d�t�T�@�}:�G�ffk� �o'�9
Q̦��ň�/[�)N�C5�D���,M���X�������70,+��?<��8��m���	���3%��w��H��b�>Q���󓛨j����Fj?�96���ֽKfZD�f���P&�uq=mT�����	
�]��X�<���A}^BNi)^�"�e��P�[5��_wg-���T�v�7
	��z���<�Dۆڿ�TC�8�Q'�7ۓ
�]�k���������p��l�p��%�����}��E�Kӗ��9���d��d��FcL��>�?��6SHNq%:�eI�J�W��\1�?�龥�Wf���e��l�\,�\�PY�s���A���
�fM7D~?X��Tq��� u�s4��(o�I^U�
����b��1B,�>m3-i�ȅ���&t�_t��A?�@��3�O#��7����^_�|nG��ƱӦ_���(&�`��c�tGP��of��ڧ���t��."$�O���ɤ���@*S������߰�\v�Au ny�H����v��ͬ�DfQQE?���=I*y��wO+`�B�I]<O9~����5�(4>�O6�l�c�:̕�?z���R��)(� 63�#π�j�����+���XlxVHYEB    1bdf     ad0J�C��.\���2@���7��
rx�������F��5�����D|�Z>��_�,�:Fp�� �����
7P#N�@?�GF�<*8�]ީK]���4�6���R'�%���cD��r�g��_r�.%�/0d���$����j3�ͪCe��&@�d4Y��഼|(b �I��82Y��]�,�u�F�й�C�G���b
�o�V�|ٛ/�V�߈�Q,�ͩ��մ�A��>䲏 ԇ�B��|2:��G�����ghj�:��(�
 ��Cd5�z��bѨ�*:�iRe��$��2Lxx�2Y)����XN���4��4������6��L�E
ڭ�+S\�R輵9^��p��ɐ�vX��	> �;�h�̭c
Ժ�	�b䳻r�*�n��]���H|�_�����Y�0�x|	� F�i�1��ߴ��JLA=�J�7�=?RX����W��S���F#��q��U�{2�����]����@,E-"`���-I���`5��xİ�yPS�v
D0x-E��u��n;���}��K���o�����`ܪ�hG:�Ƚ3�Z	՝��|ߝ|��=r��?�DU��@��ۚ2��%.�ʥ�����P�]u��b�C��,�,Rl	�W=��yE�$�(�{�9�� (f�Ƈ��>�*q�1��h|��7WO>����"��s��MY�[���W7��X����i�cn��;�B�����������'t�Iq����5O���rPY5l/�0X���rW��1��#���v�����S���@���
��QA������d��Gwb���F�}]�vNUK[5���w��9E�MD��u.Q�+�������$J��T��j�y~�מN�=y�s��z�-����<z����G�Zy��y|d/��r�����a�5ّC�9�I��~����TnR�씦Җ�gt�jh����Fwͫ��Y�uK�����6�s�����b�i�J��7���w5�/Uh�����y_�\�&;�lh��2uevt\h��B����ųr|�g45ǹF�Iz2ܓ����W&%���Aܪ$��LU���MT�
@/�\L�I�i��/������A���
ޥc�z*<�h1e���g�3�������M�zɶf�D��k�h���`!��
	5fz �%EV�!�o��o.�h�eJ�n���1a�����O�^�ɔ�3c�&=-Ǐ|����\�ueǓ�s3�I�ct��+�A�ʜ��'Wށ\�������C��	�p�g�n�������Bۈ%���l�X��K�O�h����B�?���i�8H�B֩:�=�D癿��ϕ,9��U��9���y���v2�ߕ�$HLB����kuƈ$�.L�k�&[�)M}�m^a�F��gY��&����s|I�U�dsB��	S>>��^/��R눅z���Q�0�^gޱn/A*�gc���51ܞZ�`7�
���w�+!;9]����67��<�_���FH"!Makx���a�PA�(���q6��`�k�����l;����g�n�vp�����uI�2�g��#ᇷ7����|Q���x�Ƕ���F��E����C0
<��
��h$�7fϢ��\�G.�G�.�S뎀W��\��DsI������Pm�J�)�N�G��"i�AS�	�!���<B��`D��6[���WK�x���Px�*���&9P4ZQ��M�����2r���*���s��{7α��ѽp�(�NzI	������d�$��v��J�P|S���c#�������뜞N!,V�a�Ѭ�g��o��Z�z���><%ш��a��,� |���G?虹�
s��͟����(�l�.���B�z��'�ßs��=�
1�2����wc��̧�Sd��fv=E_����k�Wj�=/A����V�%��+��."���M��ChZ��z*<�9-����TE4����#��n�J����q!
��O��<��><�*�R�g%�+>�աl?2���%�~S�U��]���|����
���E�-������g����r)�Pp�R>�`T��f�u�"�D�9:�
� �=3�W��;]�l���7k�P�NPgH!r5�����J��j�yr�NF�.�7ʾ�\ABz���<oڌD?�@����:v�-S���~�[�щjŏ�Z�H�+�����İ�_˪�
�ߌ��;a_������9���> u��Ϗj�L��:1� ��,�dh?���~��mNC��/:�e&OX%�IW���� �u���3���k�{;�����J��hׂ�R�zI�ѰQY���I��PY.[��^E2�p�J�U��P!��5ɶ��R0)��2Y &�� 
 �����u����@����@p�*�!Ga[)���l�a-�2\L�s�G]�v�pF쩿��pnc��*.d�v�8�����R=�"�P[f-}>v��# ��ދ�����F.d.=!f̛肫!,[|�>&j㌁�c-��Յ��G�c�B�.d"�½���7L�P��/�����* ��V�	�����%���o�rs�ߕ!��V8��4����d�}�Ě4���ֱ�;N���F���e���i$���!I9��2�^˴��;_
�o��7�T�1|��z���e:�z�Q8O{7dp�)�fV҄�g��EH� �֯y#�bt_�=��"c�Q>2f�8�;f��o���Y�e�%