XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�S�y��J�b�h�?�����}�[/o��;UN�&�f�6������2��Z��i�_�3��.�nY�J鿛���Y�}�t
�;�����j�B`�U���@Hr]C`��X����U�"�o$П�^,~9]�i�ϯ�TV�C��2*7�$�/�������}�,�f��0��y����̶k�K�:u)|(g��Q��=�`Hp���~� 1Nv.�ŃD�j3�]P@�K/��S�dx8�yJ�@~�rƸv�SS�j����[X=K���0�X��Oh�e���V��|��S'��i4�IB�,'KUݤ�� ��J��+:���ē޼�h#*y�+��"����M�K<b��A�B���i�`rOT?�װq�$�й���6�W�؈t1`1dqbH0��>�t~�=����B��䯻	7�I,�̴����@m�8џ�}���x���(��&d�X,����,��6(l�-η_5PЙ�H�[�	)X��F�u�@\�&\�ꍅ�:5��e�z!�@���� �t�N�}����)�qY��x%5j�#=fG<����`(L5�t��a�2uѺq�0b��E�V�U��y� O$����!6]�B���E����0��ːW0����@�*�GCI��DZ�i;�޷Z\m��q֝����/�b���tW��J�O�
���ͼ��0�A�!V���3�>ľ�*�tz�V+<!�?�"G�F:���S��C��+K�뾊Ă��kzUvR��ϱ8����C����R�XlxVHYEB    fa00    2c30�v�m���'����X�L�fB�0JFc[&,�p�W�����~�c����e��8�=�������:�L���+|��<�j�q��QU�{�|g:�Oj ��3�#�a1 C�{p�{��Ú��$�I��e͓
��W����l���zk�oW3��pF�-�~���"����� ��| �Qܰ+WZ!��i�BE*��
��k`�}�R	M��B��bnj�W�T���.��d)+f�%kN$�C �7�A?���z������kP3����3y�#�3UA��čQt�����D�T�~چ$>7gm��1/���l$��C���E��i9���`���E.z�Rz ��%ha��.S~3C7k݊tr�!T/x{�����jd���j��jj�8�M��-۱g[N�c��3�ѹ���`�1:�6�kb.����D����m�r
�^|.Q��Q~�;���nh�mF)���.�A4�
ː�w5�-^��CwC��H�����̍�җ�eSat�O���m�p��Z7��L�Yo�=,eᔽUZ�O��|C"�z����p�&J6]0��R��#9��Lkv~��LL�gf��V�_唉05��`4����/{������&��u���&��f�e*6��po��Ԣt����mF���U#2�^V	��G��W�DKت�� �X�n�Z�iļ~��ޮr�7�9��>�99y�|sTky�B*��IdGDv�)�-�<��+�Z��n/���*/� t�O�^�9$P�	��8��]<��0���#�rdÌ��JB���9qȰ{���ŭ�&F�ڭ|���"a��J�f��yl��}��	z�G�=��F\��+�ׅ��>w��^�l�LWr4�/�#�������[!asA\R{V�¸�D��
|C�����J}s�ҽ��i�Ce��	���&�#!|�ҷ����q����٨�=ǯwL�;��I^���K���˧S�#��m����~�Wf5bE~���u\5�cA�\�YL�)����ɡ�e��x�$�Y8���VeO.�b��7�`�}�hu�\���}�m����J~�ax��3�Nf��������s!�Ѕo��V�,�fG�<:>�J	�wW�B�S5��0����$����էG�w�o@b�軿.Ϋ��^/��6�V]�Q�Ĭu|
�ƻ�X��D75x�u�W����q"����Ԥ�^��<����l�(_ �q&xIK���%׃fA��Q�=gH�s<�v��n�f+�9�
�0z�v�f1�-c�6�c����{N��T�<x���������d��"������V�Q��LFĠ�B�~ ��ipF��Z1&p�&X�:c���j��@S��M:���{�~r���dU�.z�ƍbZ6���Y	��[tt�׀Ź��~ڭ��t��7���ϲ��{v�YO�3-�Д ���!�	�M8*q�v]���o#A���B�P��H4��(\�3
@����`&q�%�:����&C�m��z&���h��G`Õ��<ʢ/�
^��N�T}�~fQ��xf��FK��፺�|�;ź��HP:��Q~�u$	a]<�;HE8������8�����H�B`;���9*_z��3t�䑟,Q�O��"�n>�9��h!�^��u�8��(?\3=%n�Mac�9J �`��f�12G�z}������/N_Q+h,A���� (�T�1R!��B�xz�����J��Ϩi���Dfg~�k&����g�%��n"���)�,���bM��
fMq�]N'f�z�7�ɮ�Y��8 	r����v���;��:S�|tQ {���pٯ���Tq��Vޚ�7:|��+@Fp���>��
.�SKFaOgp�a�mB6x�:�F��Nf���I���@���ۤ�3�(��ߤS��9#�|v]A���<�����<��bH̗I�ؐN��+HL��Y�b��f_^��9�ñT���X�r�!����6*��k1)IOq�|Z��LA�0�8����4d�]�ܙ�8*�û��*�f�K���a3�b�W	(k�-k�Ro�ø�J�,��*�>n1[4j���j6\���s�}�����)�]&JgDɞ�̆���0Uv��v
�JWӗ�ie��Ky��]<�FL��ߜ��ç��@a��:տp��0,���|�t�{�D�}qN�}g���
�z�*�c��,������9�lA`U� ������C�<�Fy!O�u$�����?w�;M���`ף�(���7��E��4��ڟy,_^ی����A@�b�pɒ�H��-]*m	��%"{�'Vf$�r�lP��!���І��_���I���0 �~j�4���aԓG~�Z�V
o5vj&।C�;���\���������4અ�:����mE����wT���7�yNP��B�,���������q�v�M�+��6�j�%����4el��=��q �羽�u
Ɯʊb�#��/���n�aiյ����͐�
a������6ʴ�tr|'�D_�?�Ɯ�w�#uu;�7�t�>H�'Hq�J(3��`Q���
ɋ��0yVĳ�Yq���� ��P��A�i��.�B��B���?��K�+N��B��/��
�~����q��R`!癱7��f���<�Lk�$�&!Y�{��!P.Ӗ�k}�����V�,�T�)\+q_޺�aCzʽ�����r���� �@��pj��Rg�_��7������պ���K1B��__��N�P��uO��?F�ܬ�O��B�`�g�F��+����;�ў_���b�
���c��}f�c-�"�̀�PZ�0�oM���q�:�h��q��sZ5I!�֎�
ķ����Fe ��2��D1�P�ߔ�V��hM�I)�z,)%%;�+!�b��i�p\\�['�3��K+Q�f���{�*��U6�6A^1Ж{�WnY�@E�'^vC+ g��i-D��o(��fc4��
��Nh� ��{�b�'���xT�z��N�~��For�N�z��a�0�d�A�B~P�'��Fl����ӑy'G�'�M�W��B��{�-w�%6J��j�FW.}!lNF(��TR6�7����L�tm����eFk���U����o?���,1$F0�j���Ĕa[�������}TL6��ć��mo\��-�JZ��v�m�� S�1*�s�#�s���c���0}�H�����!�T�F1'=�(�١d�G���~�N릚��W��W�YH�/���d��0��gaOH�_sǓ�,�&yK��6q�SvB�hU"vj�#)�=B8�r�j�_�Ԧ���m�78�ǝjk�Z��>��[�? �v3DӟHd`qA�(�R
J@}?����#6Zt�đV����#��s���*~�6í�)O&t�+:�i�ۇ�����R<�f�!t�sD1b����������DT�2A�|G<:2?��'Q���W� �Ig/�Yu'\��z�2��`�m,����5�4���<w��;�8
y�z�F���l�3m�t�η}��r�r��h��;��x�Ia�_����JZ����������'�H������*�����pV.2��0�(���U0��\�gϗ�0���Z�h��)��߮�͔+�-���>G��U�IDp�,f#(M��`2v�h	�!�n�L�y�H�mS�#/���Z�L��f��wW���ѭ�4��0I�q��B��i��-�ș��PrTF�?��K7I���e�)��R����n���!C����ۏ��ñO��x4��H��a�e��z���m��F�w��l��*��������,���ĊG4�;{:w䑭��q���K<��𴎦��G�.�.ݑR�So�����U�����o�#���A*�mJZHlU::�m�z�?�= �	��;�Q�ҭL$�5�q��F&�0��$���s��s��$x-a�#P�XC}
˷�jT��[,SUr��|�ұУq�A]%*NOC���A�v��Ə(�A�贫���~ܚv�z}�z�&:�`)O�=J��%���0P�'�j��#��7�q�Y�0���9c%�u4]M�M���TM��>E�O�_%�A�h��r�!�<^�u��}3Q��C��(:���J�z
�����153�Hc��K���yn��ϳ����A�&|E�Kw�p	n�,�,�Sx����H�`�he�r��O}v���"�����_�{���J���<4z"&Dw'A)�����j�l���\Yx<ʋ@T�?�(��_B�n�ڭ�����6���/���q>�+�p�I�E�D�	r����S�p�0�i�t�<����n�\��f��]jӕ�オ��iW��34�,��3�o�U�/�$�S/�Aq�̬� !�L½�mI:�U5lB�87�;ɜ��^�('1�ڮ��~���?�٨����یbۉ���
��P��ρЇ�.�%�j�#�C_I�6D��@�9�������<Yh�g���(H6~�
U��U'��H�2�K���pp�P� ��;`�׶�̠{��� �6����{�OG�~�gFSt_DQ:�l\�M��'�'���;&I���������=ȓ3Z/���lE1��w��>cig�ڐt��"gm��ۋ�4�	�tisGAk9@��L�/�*�I^�F+T�q��E��sr!�Ö��8H#�#p�6<k)9�O~�q,��1}���?z�|��]mĦ;�[ �0�m��~n����Q �����i[K�K��=�Jn�6� �Ƈ�S]�"�ۊN�u��]����|�]��i�����<?[�'�Ǔe���~Ǫ�$����#{J2�A��)tߑT��C6z�YX�`�a _U�v�!7�9)|��h�m�]X�����'_'�a�f0zV2j�-����
���V0��/�>�Q/�@��5 ��Q�	"3%'|������6s��Ƞ���9k������}3D�4��V6�v�IAUK���I솨f��r%�3P�jH+����:�PPA��/k �(�U��uK��M"��U}��z���
u��<�@�g[���X�MV��2Ng5d?6cN��	��������*�y-+<�����z&g�qb��y���Ǖh�b$VO��ʀ�m���i� �
�&c��( �{�(e� 2�Z���[ּLf���F:��^boΜ��B����y�Ol3�l/�;�<׵[�B�;�A �[��\�ڦ�M���:�aR$�'	�h?���W�Ilx�������y�f1�V�J/�2�+b��lB�>cO�������ͬXs�y}<$%0���,��h(w4�5�`]k��`]h_$%3�S��?�o���w`��{�ןfĖ=�
�u���Ύ�M<0�i���0�ۛ�ib������2)�b"�o�x},�M{7�8�ӎ�Y�V��i���x��(��f��u�URDy�c�9;��R���M��4=�oUf��K3����Ǣ�8��h�o]wB.q]��=�0K��$\�O���{bD�@f#[i�z�C�2J��p�Lb�&#�y8'd�]��2�NR��Q͊��c�:�� 	��]�J��i��|���Wcl8�W�8U�]*��9�/�:h^8�r1R�[&�*�=t
��}�Pg�m�S�	���u�{4��&�!�����o5�+@e����a+�g:�T��9a����h�d�6�;$�ж(U�y��I��:Y5�E����[�������D��3��:��E����nUKS����z[mae�� ;�Hՠ���V5�o�3�LN����8+ŗ2T�*?�v�?6���[?;�xj�f�)�!;����>���;� Zq��l�n���|`?���K�tC��,��d?
�_Ψ���+o2����;T0�EgG�UU`J�ȨӪ*�v<~/����~�QhF{�[m�m�l�r]n_�?�s�iM>�&�xf���^n��Vt'��Ƶ'�9W ��;<�����s� ,sG������-�������a�T�j��}I�5n�G�3�L�m��I#��m+�~�5�Ơ8��6~o��m�BH0�����z��D��bd,���U�kk%xeFuڸ9�P�p/Tk�<������;���G�\\���Z���2�P����X�vl�����\A��Na�F&�$�Fh@rX��ط�Yx�P��� m��0�����j����s��Vc�U���&�;Ɉξ�����;��ý����V��mp�PY�__�3x|]vݥ�ٻ�%���"O�=WP�i`��JR�(
�ID ���.r���S����Mw��q$����$���q7���t %��R�I����t�R�bxY�U��.���k�KW�se��+h$A*�tH�,���-��auQ�.~_�N����t�#,0%kc].Ɣl��#x�1��wXx#��`	H��Хtg.�߂��pV޴ 0��ѣyz����	ʠ�v	#f}��d4Y9���Lԇԧ�[�)3����ps�Ѻ⍩�٘P�hK��^��8Rؖ���(��÷�i)��ӏЀ�"�"��}&q��|0s~�q���4�'�����<Tl��o(濭ۋ<U�OC��N��}'�0~����5�X	Zpd'*��\i�6rE��Oƅ;���-�����"�0�	�i���tFT�w��r]Y���(L�N����5D�+�ϟ��{�^;���ߔ�Ц���:WʣT0�����A��7�df�e�
#��j���Go�O�4���ܡ���:T�dV�W9�m	N��z(�Z�߯�g���;�Os]�۰<�z�j���8`<���#�ށ��&�}_��E��/��U�c�?�>�
�K~oP �q��#7����B��໱9�Kf�L�T*,�UB�>�㽯w�ᗔ���}�L���N4V�� GY� �4�\��څ��E���L����Z�K�-�)�8R��PGө���֙�4��������g³hR�=|��Z���(�̡E��t��/f^q�Zڒ��MSz8�W��*/^�� aH�����{��w�۰��YM����h�w;�Ÿ�0���[��#�f��2I
�K�r�Yd>���{2�2�ɓ�F���s�jQ{µ�ʅ����c�]h�)D�Õ`�W+X�x���ݺ+x����DA
�WB�}yK�6m#�ܞ�	2��ȝsc4��)Mv1,�{Y#�X� �v� \��pP��}8�ڪ���;?"�P��e~3ޔ_R*�1�؋|Al�<�cd3u�Ԛ�@��&ܨ�>7�4���ῖ���ˍ�Tz���flx�a�[E����>�*���u�5�edBq��n�e���u���#�F�t��y�c ���]/[⚵��8�b0���I&�n�Ʒ�s��ć�猘�L�ڄ������T�q�r$�ʿ7�?ȫ�C�� Iո��x~�\m��s	�!V;c��������ߔ�Ayx���z`z�2���5��FY�2�=��H�BQ7��~�@V�z*7��>߫��>̗(�Q9<��<��I�� ����d�s�s,v��]4���<��_��:�]��\��V�M~�Xl2�;Nࠌϼ%� 5����d-k�����x2�|�HR!ɲ	o���B�+�-d�aŝ*11-�A��0Q�x~i��e<vP�4AZ?��6�( �.�8�^
o���a/�_������l�C�H��u� �p-\�Mq��M"{sp� ���%B�D)9(�Q���l�E@���N+�W�&ImQi[ؔ��Qw�� ���8J�w�L��xNG�u��+݊�[e��|�l]zT��M�d�0����s�\ê����T�#��}&c⧻Gt�2���&l�eȾ1����ѵnY;`��� UT���.; �#&����Vi��uG���C����:��4u��ƀ��w�~����ƪG|�hyO�o����cT����.�����Xd�q3���ba;�2�mdH�g�e���wUa9SQ�]b]�IF�����X�a��Tٍ;����0��]I��\4�P^~�#�K��u��`6]"�>����|ٺ]�t��sM��Y�\���F"~uB	k������ь��I�3�ݔ�F�U��P��֒N|�,�^����ʃ�(�<���?F��{�T��d�
	y�}�^��g�0����k���{�x�J�<�p�?����E�9�V>���p�J�0��hU�<ɬ�=κ��z�Q	�0_VY=�t��4�mE��'��𑆪$�
�Ɖ�|�U���	!p�'b���`�Оҏz���P��Z�М�6�5��������y�!1Ry���r��}�rs�\x>�N�����ZГ��S�M"<��I������cgu�"�q�;rlIHT���b߅��g�+�۠
桩E^\��OH6UqZow�?��w�Z
5��h�u9c�"�6�t���ˋ�4�`�R�;�`��I��$4�\�Q��MиR���/_q\;]��?�6���Q�0m�}0x$*L��K)Q}�k�4� ���0��x�3�U1-C-��ν�m۶�o�S���~�Q?�'1[��PDw�U���	�0?�'Pҝ ����lp���Uet{\��E^z��	�U'��M^e�2�J�z��a�uB����4��&�����dCv��2f�ZMW��2X2����.��Cr��G �c֠�mC���D���r��������?�W,�q�	�[�b���!�=ݟ�9�U�sn8�r]��u���/a��k��&���'��L���P��RȾ緇{��k�����٦�9LiQ�K^��[���)%��=C6�	��p{�6�T0c��C��ՙ���(٪t+p�w������	��QGf9��J�S�o���l=]3��F���͝��X�bϸC������R
�X�%|M�hL+�>�̫�uվ�9��ʹ�_OQ�4��bx�տ����'_�~�K��:lI�����wGw$
F���C� (��yPB%bK(���c�>���(���y�c(C%�.��tU�N㻩(wk��~ �pH�g]uK�jԿ������ ���|5ăP�t�<P��+����ܧ^(W[I�*�������X�o�=�G��V�iB�>��Po>	6Ѓ��d�J��*��Ɓ�j�,��TRwR�=���ߎ؅�H����Tb�B�C�%��#��#�TD��Ca�;�#W4ii�&� x1�W���@5Wܗ��e���s�:1�������_ W� L�Q�=؛�9�O�#��Y�Dj��Y�pR%=���F~u���
�lT>�S�#����a�a8i�+<yA}��*S��"�ysM�� �0��&Th]�j(���OY����f=��D���(���O�$��r�D7�_�#�� ��/aaf�`��A#�^e��*u}���Cv�JE@v�=jWJ���F��YS�(�ouwHAH�
 \P��S���A��Ꚋ����=c�FCV�h����4�;Z���q���ֶ@1Z%�+�@`��g`�<�B�8�J`��^���K!}�2R ���&"��|[?�z��?9ȕe���[�K%��U�p�$c n��U#���0t7-䡏ezsAW��\�[D%�T7��}���t[LN��Li?yq: ���2���FՊF��*�Y�l�H,�U_r5S$��:l$�G6�b8%v-̡i81������N�-Wuȑ<v,8r��ۨ�b�e
�L=������|��Yu۲�1d4� �:g�67��@P4H]�x�� ~��j5#8����"��f��'s��S]���vt������t����i�2l{I��Ǿ�N��8��62��l�I�D��y�ztϢj)'�Da��V
��Fe��x?Qj������S�[�P7]Ẍ�Di�%2(#g��7�eNb��^��m���l�x0�z������3p����"cP/P���i�t�Π7~Y�(�~x�1E�C��ȑ�B��잕�G�w� ���d˥b��$_�z*��S�^�{�0��{���H�\p��'*tV��:/�ʼ��d��2��R�.s��N�,�F��M?��9q�|��6����`����JZ@�u,��߇�C�x����H�$�j� Qԝ7��[~��44������ǝ��]�H�DGkGz'0������'.���;����ح��u��/�@2߬�e甙�d "P�(���ꞙeĜ�.l�K�[ Wѫ�#<�ȅ�\�.�6~dYD�$���0�6��oZW'Lj��."���v��V:3����`�����9t��=�Q�UP�:�J�Qd��f����!2�[������qO �3��Ⱥ��;����8܉:��xwjƍ�S�b�=�g =D�V_q���mE���2p����<ױ��D�$�����x����Tp��rκ��bV�6�2�����K���w�������靹�%����{ҩ�5�a*M9y�,��U��'��~��[��S�$}��{!�$��!�ᩄ?m���>������D����� ��5��CZ������+�j[ܸ�B/��7��9�O1�L�f7ʳ��p����0D�
i}��6?�&�;�l�"�	NQ����l �:1�q�#5��0�} �&��6�;�(˂W��<j���^�͋IS���������f}/��}W�,���:b�}�§a�rmԚ(���q&�{@�4����4 �l��r��TU�'�L����۔>g@(Ul�����z>�#A�aGNFf���ݤ�7��	^5fw��썅пUr�]�Ŭ٬��V漎�*J򔞵�\-��Z��.n�������nG�3�zw��Ik��7ܽ��K�q|�>�$D5�o�<�{G<熬G�Թjp�Є�)?�>a-��Ae.(��٘U���{yǑ<#�O�V&�N"��}���`�x�f��^l�;+l������i `�H��O��^q�b8�kE��N�n����>$qDt�%t8�%�#�x уiQ�<O3������Fyj䊜��2�f����3��5~:a��B�L�@S���Y?P.��?{)��?t��4�p]	a�6�!(���\����71C�
�.\~���n�E�� �gb< c~%��A��U�[�4�~ �ɔiPU�Z�K?��O����	]�\mh��XlxVHYEB    1e8c     710ui�Jd_ �@��Ec����u��U�p��O���ʽ��3u�U{~���Wbw=��h\
HҒ��Yƻ��(�RÆ��Q����&�?
5����u8I^���=��*JJ`-�h�k�I�tP��aq�X2�`_
s�W�O��Ũ���}*�/"rE�+J{��-5I�!-�!�^��2�Q�ϯ��IXBJv[�����f��%�Z�"��D�1Ol��h�W%�E.��x|=o��B�/r�lH���w�7Te�!ɀ��Uk g�fd�	��ƽч{kȥ֒�9o�/������jZ��o�}�,8ߚ��̫2c�����V������� �(`��w�y�Y���`��\54#����.�a���?��g��dP��V�lQ.�o�K z&,�V���:�UM�vC��Y/)�^þ�����r�tk��p�-�º���R:�6#������m�Q�.8b��Q�6snY���U>��͈Y���#�p5���[�ǌ���ev�W�3�5f���\�[�2R@`�(^�Y�lo�P�~oH�G%P{C�����Ac����k�+��U,���oD�nʜ_�L����Һ��(%%�#/��f���q�313��3ҷ�x�%9=G␨��&��G1�e2�iU~e~��sS.sTh��h�EY���5Oc�&&�X�����/~T�8,����XÔƳ���sф�^�'E�� h/u��O��L�mU�����إ��z�^��!H�*�dT�Oi��T�����P%���]��W�����Kx��e^?�檊�	�ټʬC!BC�Px<`�1,Ek�#�k9�Y%|֓�����^�� ���~�������pn��:Y	���@�X Q�-E��]h�Ml��{�K�Pn�vw�����E=� ��d΋�?�&Ep(}����D&|�w�%�Lv��f�ԡ���2�o���)a/�s�_y��+9��3�0���=�]��t�AD9:��#�t�m�I���}�Y8��l�7����7j<ΥA�r��ӯ�=���/~�OU�3��d���Z�s�F�sU�ִ)� D�)��Z��� ��x���s<�ƒwXt�������eK��C��r;ʎ����I�����p����f��I��ʏ�0�d4�3�s�]ؾх�dJQ#sc�ja�QF2@ V[��9����4F����̫���I��{�VVH�p&��� �y�E�Gğ�\��o��>G��]�xL���6Đ&:�֌`=e����=rT�e�r,���l�Fz���׻��qS)���k��5:T��43��*����lQ풱��uX:c�6N-�pd!�R���b}�@�rL��UY�<�2�	�1���	�H�k�����p��4x�T�}�	���+,7�'���Ё2�S.�:� ƻy�b!	����b��S��DG
���U�Rx}����Ъ���N��m��h�ė�v<"����O(�W�.��n��f��,2����"�T��Z��Av�?ˎ�����s:+y�RGGHԧLg��^��'���������� (�����������d�Qvq_B�}]9;;�N�d�9��(�;2O?�K7���X��t~&�X
ۣ&] #'�[I.���������c�&Am|=��wK�o��s�#]�r�T> y��n��ɤ܊I��1HI���~���p���[~��sp�N�6�4]/�I-|�����U����yG�^�r;��J��2��&�[�l�1c� ݮC^e)��@�<��	�Q��\�(�q�F�