XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������^�Gf���2�!e�h�Q�
(oMd"�����I[�[RC.��d-����s�B��#L7�g�A!�a�Ñ$�2t�g}'�v��kFɕ����s��JΕUߌ���ȉ`OX&��ר*j��	&�p��O��ms#q;�t��7ʾ�t����e AO�ۈ��[Z��o1�ӫ�v/�5�{����%�M�S���*�%�1�=�<��N�[2�b��A���ؕ�������[U�3����N��8���l�(��n�t��Q���b[L��Qd�t�����|o2rMN������|s1擳��;#Z��P��@���o�0C�x0�$X��9�X�:�GN�����>��R;)!Tt���<gӁ�nu
:An�\[,��K`D��'�L�6� �#�>H-�]�ʺ��.��s_����(��b=Qu���p5��-L@H�I�`/�� ����u�P���C�f]�u�"e�	v<�y�q�.���O�>�g�(�t�x#�HG����	�^�0m�$�n��~�(��+K��C;G�1I�Z����k�Χ~�I��칉.K��*n��"i�
�.�!
�4X��lV����p�d��
p��a�DdE��Z�ޢ"�|!#p�=��Q.)�a�����<��D�����A|ga����1��̯ �C Doh�y%d@���'�_;�����)�,5*��Z�)���$�H�ܦ(�|�^�D�(d]�z|Vo��-�N�ċ7D���կ�^J%5�ޟXlxVHYEB     872     290�_[���Y�B��Km0�X/[ЄW2Ϟk�^�4Ӷ3�MF�/���nt�}�ȇ�X�\m�Ԓ��"э���s�c��s�r<��e�9�i�oST1f���"7{�zΊ��騪��K[M�� C�d���z�굠�9����r�m�a>�w�	��c;���{�\yjH�\�]���~�U&��Ɔ�h@��0R����h:Ǘ��:v=?��l;��*bƶ�㋜�Ô 4\!����~9����¨x�~s��a�F��X�.(����N�X;��ۖswT�d�_�šXl�>�r�"a][@� [��Il��T�yM�)�b��f/���!�i;S�Ϳ{�D^��X����4���\I����@}gI�4vL�h�$��tVH<V���OJ�P��g�EA�Yk?�
A���y&.��S���vYuJ!3[�n���
K:��+���n9����J�k��w��nel=¡�s�;���
�Omjܨ%�;��TJ�F��)2Z�]�:�AV���O����í<V��߃M�#��� �C+�Q5\�
��70KLDH�}(FT����AXlE�
9(� CcƁ�0k��>�5��x���F�p�^�K����ML�/�$�B�����U�q�TЏI\���Ɂs)�U{�&5+��}�"�2O