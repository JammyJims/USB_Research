XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=�-�,�/��m)^4�a�l��Ƥ���O͔,˃rrf('v�)϶v�n�n����;+��"p���i��k�����5�H�쬐����꾭�h]�l�*ȳ��iy���]B��V�[DZF�{��L�\�����!9��n	��#tW2���t@���+����5��:hq�ׁs�](^��� ��%�~?c���O��c�K�O��,�A��X��.���O����"�����gp�Br�����-���:�јl">��j�-P��b�X/8���1�!%�sb�h�ct���F��l����y�g7�OՋ������1��L�������DS���ؾߠ�T���hr�h���co�=26}�3�]ꍗ��<a2{U���B/���6�r��-p𰼫���/(�h5ZcM��c����	����;�ҿHӑƛ�0�I,E�7�4��H)J��g;S�v�C_�8Ƈ~-3>��+�,X��Tr;2ϥ��Yb���i�#��<��Z�S�bb���� )'�3K����E��2�\F�b�a�94�Xl�`�r1X��j�5.��Ɓ�9yO���:%Yj ���^�9���Y=YQy���)Ԡ��B��?,��ʘT�h�}c*���!D�&� {V/��d������{ƕ�.���� Oo�Tmm{b�w ��7�^�i�I$��\�㟏�M��><�4���;�,wc.��?=ˈ�VVI�b--a�!�p�~(��7��+���+LeXlxVHYEB    25bc     bf0G���S��V�|V�3&4�\��-��PF�Xc�%F��*���p�ә��"c�����8�֑_�ˁ�����0��6�Bt�'�B�_K�emdb	:��8P����L�NIDI��(J���ʤ��ز�TZ���ͮ��ƿĩ,��=���%O�1����8�ea�91V�Sw���c�a
�+}f5����5��A�9+(���Ǧ؄�?aJCI9����Ha͔��g�F��';GO�8vU{�P���J�t-�S>c��?>77'
 @ҫ2Mnf9�8O��l(;���=�<l��.���M�"���w�Dr�]��ED`��r���_�Ɋ��V��͉��|�P+z��p���^k����U}����E��F�sR��奄R�fծ�!��C/�OP�X 1���&ރ��a�&�O��%|�A��g���*�z��^W,5��ٵ]�HR]����p�����*�B쨚�C��&Oi�MĨJԤ��&tY��K���w���}!v��B��Zdn#͋������h���%�pYW[��5�Z�?^K���}�^�y�}� X����|͝)��?ҧS� 6;#N>��n,���AG'�
�m��WOgf�X�G��n𥎀��$�C�,2�yB��*j�/�\
9-������Ŕ���櫥���]��� �
�����XY�Th���o٥Z�޲5m��8,�]r/ۈr�Xge�u"8e|��}����W�KX	�N.p���p����q,g�r�.�@[��[ָd���Y��f�������ެ��g	m�$���!�L������v{c��( Z�0��G�ǡ�xc
v[�35$��:����,�h���SU������i��ߙ�
�?�{35MinA�{�M!S���/�;צ��3�0���֠���u~�T�P?k�\�s�H[IhHCV��<��5)$����Mnp��sʑKL�h9�M��M���b�����Ю��kM5��T6M��[��I�;���^$����d�����1"f�}��1i�a�����^e��n�%RG,_�A�Nn4�3s�T̖�'�:�fj��m�L��X5�z��|�V�]T�"�#
ۓ�w)�����y���H�xLUA^�ѕ~´(2R��Nd��E@x8��	�ݪ�.�MzI���=u����5�4�8��^�>ѡ X܎��e��5�-�9���\��n�'#���Q���`~:�$��"�rY�� %fպ�^�4hk+6��6��;O��\Fn�t7^n�Œ�3�Nv:T��P�)ۥ�}/1�8i|�Y͸O�bM�Kw�>ըx���KK���}�΁���Jw��jk�E�@�FQ�c�謔�!�r ��K�ŕ�>���(�X#�d��+'�#�y9۵��n��.1�Pްr�!'��g�K�L����i�N̆����g���4�8�S�!�[+�u䄹q5ݳvٗ��Fp��� ��m�}Z�'�C��3����8P$}7������m�,�Ǜ���=��s��+��r�h_�׵�g��K0q�쑵�.�<��z0��O85=L^*XM�ti�G O~�/���M��|��k��Vd���5������SOBqׄ�Z�͋з�O���.����
����?1V����C��tη�!�y�:���ACz�	@i��z\tFMiw�z �X�w�5X~�<[�i����;��_ 	�ö�/��P��}�rֶ$H�Ҽ�.�fH
[�_��(b��M_ТC�`����v(>f�Ƙ"[�*��A���N'׾��突��Hu���~5�� m�f�`=�#듐]�IP���p!�8wmW�����kJ0g��c_[�&t��u�m�Zz����*��W qkf	I���:h�_¼8݃�-��!S��Ap��zS9�m;���_�/�H�D�ϖ�U�c2Q��"������vaٶ��_��(����Rd��"K���y�f��Y�s���~|�C�b���Q�IF���A�M���[˗���RغE";���dg!L�>��a�P]��ML@9�jX�v/|<��ۘ]M��Ӛ��C�c����na�/u07#���C�0%�o/4f�g�ӭ��[{���J�%��]4�x~s��x�
j�����8��ش��%f����x/+y�ќJ�Zͮ����OUS�LX:VH�Nbj�D���qz��Ω��Н :��D~z�B���"'#9�<;�r��_ �����\�7�<Dx7�o�?�;[��77�v��͊h��g�E��BE�98
,.��H��""�X/D@k�� !ǌc�m��-��3���`�_{���p��XO`eE��Q�1Zz�`~s�Gn\�J�b���>��s�cY< ��]_"�(���Hě�9���G��Fc�+i�c�=)g�^y.INf�(FS�)����辞m6����&)E���|.��o�b4�b�.�1J�yOנ��M�6Kd�S��x���)#��U�HNuGw������!��7�7�TR���2.r��[�	��CYg�����E�L�~�G#rW����G-�+��g�nJ���Ȩ���]Wa��_@	/���w����k�e�oO��Ҹ�|�Z8]�?Y����Z�͚5;"e)�G�;D�Y%d!��U~1q$�I��/#�G]YF予���(�S���%-H�3>�v`�`M6Th�O�t���-j�@���L��A]$�e�,�f�7�nyP
���yڛ�P�䥗�Knr`D����y�_�ؠ�ڛ.}tio�	\/���)��Rb�u��)��F������t�ΖeW�CY��?�c�.ܓi�����i�JMM�}r�Q�k�����:��^<ƍ�ѐ�����?���(Q�Ӟ�V�bh��;vrS������P���H!��od�D^��!c)���o���#���^L�Z��c�%�V���axK�G9{�A$��K����7�g*����?h� �E��
=bcT� N�8�'���i�@Y�6��%���������