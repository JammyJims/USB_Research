XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C��;D�n90���"�.���n���#�*���W��Pb��5��vhWᷥ�x�y�O�6�$��������w�D�E��]��QڣKf!�w�M�TK6��6L�K�{'#:���^��\�q:���v��$��P�����t���d�hy��Y����n.�r�&�^�J1�]�$-����4N�����U<a7��bD#�؏&@
�D�SӰ�f��E�#��KQ������ ��H]���i���"�ա��-#>|����(���>���{��E����Hd8}s�Vb��#�p�m"�� 
RL4jQNu���pΌD�A�	�M"%C~�Y�XKB[/�� h��,����Vcpq���W�~���g�3a���l�#�ug��8zlP��}Y���ؙrH����D'�f����f�h�C�'H�!5I>�y���8%�d�kN��͉���d��=�CVcZ��k��/M������oJR��P�Հ��<��h nף��y���Q�4m�TZ��]�/l6�;��X��|���ߩ�xC��9Sd�.TM%�o2%S!R7�GZnn�>�G��zғ@���mqƑñE�a ���o���(�g+�ix�lz<x�#w��yϷ�`�b-:T_���_,�?�6�U�M�Wݔk)lT�{��:�#>����������`�C�4H��4Cl:σT#�����vN���[6��ӵ�jB^��T�o]�!�|楽��WPHϙG͙�%&FV����24XlxVHYEB    da51    31c0�k�$7R�΅����]�����Ԫ݄:������AM���>}||��k��΅����.A�6��yU�7��>�>������#�l��!Ԡ+�� 8�w�u��m�N#�X�d]>ߐu������R��Y�V�S�;�ҡ���d�̖��еЇ���^�2^��Ҝ
��C���4%<k�͕�\�a}���}AmU0z�҂��PXT߀,����!$EzE]��d;��.��f����Hx��s�-yQ���%?��ī#��<!l k?���$���6$�]���~wS���(��*y�BTZ�X�x2�Aw{X���97�b H�V��~u�eqo�
�c,�Yk<���؜�����$��!-%
�|�ܴ�A��,�r�_
�Q�ݩ���֘Ќ΁M�hl��#�PG<��D�և���˅�$�R���ᬧ�n��K�9�Aj�ّE<����m��uE�W��BU�H��ن\*]]���_+�,��D��t�;~�@�mӱ���|��K�	{H��o�%�i���Pg���5���Y�R"h��ZDl�����[��� ��SP�|��oР#qo<�S�ӥ��]PA��U[��E��Mn��r�������Ms��;Г��NP^P����Ĺ@���	~��h�_j���m,����"�<֚�L� t|i6+��(@h��q�ٲ��*�l�y��:(���3�u�P3[7����;��ʔ��J�
	nއ�Q����B`y�u�l�.}7�ꀟ���9��Y�WH��?,Y	[�}�%�R1?y9��m��vn�XX�x	��������F�cj��WNE�o\��	)�9���LF��ܨ�לd[�@����k�2�)���� ��yDR�S({�R"��VpHl~ɰ�>��C��a�ͣ��N���<���*Cr�u=���W�0W����n��Y����y�n�X�Mt(@�([�y)Lm�v�m����:ټ'60;HWM;Fn �.7R�q�	��:�!�2*�et.��.�\��^���m�`W�YwB�%���$>�o=k���) ��Ф^L����)�����e[��mk��p�^|��,C�������A?�o�������ygS��&�N,�ǿ��nˋ)���hD�n��?�����F����M�4��G
��-b|�rx�{��#���M���x�h�-�B��͑d���C��
r�U
�F���>a�eM�a�uV�6.�l!j �J0+��yV���!���x䉫=9����v}����!��_�瘋�߇��{w�S�'����e�������"-�օ%�e��q<N�[��P��pdZ��Yȳ����4<�(���4�˕x�� ��� V� Rq�(#+RbT; �߾@���B�����4O��h�$	.�� �ch>7&`�zV-x#3��U���5�èN�Ү6$L�]ƹ�}t���O�=(�\�eY�A���s@�6L`	�F���ka~a~^��:&�Ƶ�� }����3��yUl̀���	7�\��It$/Q���A��1���l*71Th�ܵ��h͜?烲��C�����.z$xzOH�7%�oPߥ�*.�W��TgO:��1�ޟ*[���x�p�d%� ]OI8���-F�s�.s��l}0��N����Cx�>����3�P�<�hB(Xf��:g�I�J!�ֆ�<lxٽ�zdϱ�i�������?�Q͆�W$��J�����A}@@k����m��)�������=]�l��ox�q��b���Qrr���CHBZfǘU�Ӟd�9��?�:���1S[�ۧ�w�-�|�#X����2��jo��$�1��,w��ZLМ"�3� �^�����$�KӀ�JvI��?H j��������i�xqK�@�����E��v��AHs-�8u	n�f��\J:�Gt��p��Zx�=`����a��)� �)k*9��\����RF��s6���!�H��%S�@db�����c�r�v�t�Q�����-��(_��1ѩ,��=����ϋ���+�� V|��������}*ě��ߨF�B>�����z��p��0�"z����1���DU��z-i���>y��}񛃃?Ϥ���]�����6�4/��y�7��^��g�|�z������H�Y0�_Ht��՞���w�kM�C�����@�J$���s`[���l+�$I'y�YP5�@�����j��sK*���u�x!�2߻rd����<�a����,[��)��A�ko1f�mU#��d�7���=�<5���5��}E.Yo%��m�j�@�!H�3g/b��|h��|Y�N�|G�������wݰZ�W_���V3�	�;]k��o
 3�H1����V����Z@$b����_��1_�%(�eu�5z���0bڀ��i����R�.R���wNF��_h�;���ٹ��1ذZz�E��#�<X؍"`W��RDT�SN4l޺�Z>R��xh�?�P��6��&�L@���{[�W
Ek��`(�� ��&}1B�L��6�.����n��քc�,�6�R��?��%�<�+��U7��Q_{���}�3�0�I \|D�$~KڒX�����)+ M�I�=�~�#F���������z9��A�P@�-�|A�d�����c���AU�p�@��J�Gy��]I�8��n� �I�m�iLm8�b�~bToFe>�y���1Z�-m!#J�$K�N̊�5�#�hx�|?(C�!���b�i/c�PK<��e�·tL;��k�k���Lc#I���	!"!��%����s�F��b̑�L�aQB�0Lz��@;�q�rѬ,��Z�Mc�;�`9�����n�RW.R��MA�7o�C�V�
�W���+�8f��T�P��8�٠AVC�޵�ci���2;� �@#=��y��6*��ߣ|�ʎ���X��N�@x��45*�Ό�̀�a\A�\JyK!�9X�ڨ&����H����w���!����.n<���"4P&����تyup6� ��A� W<ܙ�U���A���dd�s��ޓ�	�xBQ�b��~[�
C�ڵ�����1�0k%�ø��'8d�/i^IO�j�8�����h���CTsݬ>
�B�R����z���L���0��T�}�"�?�鐏;��Bl�� ��{#ϔ�:���4�1�Z�M.Vo���@�m�^�&���[*��B�f�Պ�	<��nn��٭���h��S%.Mq��T�}FE�?���*x���0�!k��c8����O����_Tʣ������J{�oԵ��04\�ז�>� @�J+oF�U���3N��z�a�+����|S�S�`4�IX�{�F��jO#�N~���vۏ*�s�ЮWd�"���Ǩ���W�|Q yc�/���(��f� +Ew`w���0�� �`�r�4`G��H��KVw���D�_��׽��<�^	 $���z�>r�q����^i~ ��
3B��k����}{�D�li"�S�Y�uC[�H��H����5�r#%K�	������縚vB�Y�%4�+L�=���sU�)��l1'�o��#�_�ҡ�r��a��5�v~�GV&X˅�`U�3��@I��F��,��0S��4YlhH{��1@_�k��*k��`�9�	��!���=<7�_�5�!��n�Y���O�a=^q�ؓ��,����b���G�+kN�!@�P�Z���#[�7�k�n9 �:XA�兡eI+Poj2MS���Z��;1�1�b�p�׀t�z��r%���DW��w{�%1h|��;\4J���o�í]{$��-ݡA���w��S-��ָ��_笒^M�ęXd
-;ཱྀo��0zD��\l�\�����Pf�cf�4T��JD62������n�?�&D�&�F��EU^)��J}�Lv)rx��F�}��>/�!o������ٷ����� �ڊ��o��F�o[��� Az
#@�msl���S/FNXl��[@�	�~� �&�i��j6�Vě�!����ؐ��-)�?_��e��V�e+��sc�{���D�-�ŕ:������P���˲���t�@��m	(��|�zo�]�<��[�[lmE�T#ad��$ α��c��#��6.X �г�>���-���Fҩ�0��8o��^�}ÿj{��/٪�7Ӷ�TE��9���֟k��+H)@�V�<��ňLC��<�Sr�20� ޜ�e�ͭ��bvM���f4sˠ
6k�l�=
�J���x8F��,> �c�G3 |x�����`L9���>��]/�CM�=a���w2 ޔ$�iPHL��)�Dm�f��bϢ�����Z��{c�v�i�ƹ�P$��W����'��,ea������ۛ�|t\���|��M��\?,1�b�B�z�s��S�s ��/�@I�k-i�Ř�NQ���%�}��]�Y*8B�O�4)�V=�$iOf�3pI^T���T��-l�G�W��T��]J#�� ��d��&���w{2������@+i�]�W�1��59�t�\a�>@��1S�$�{�E4��r����q�V+6.�DCQa�蛁	)[��t�w([�^A�4.�@��gI��ԓwFS���}����S%"�B!ُ@)�b��K�KSr�h;��3���&U�z�.˼k�Tw�����|	��ÞVWq�g+�omC���I�hAz�o�# ��'<Zu���O��峍0�H<P����.A�X���	c�To��WT�mC��t��;{b2z���c���:`����A�M]�&���cq�$2�)މJ'a��g�m�,�]�V<)Db^JW��hGl��Wg*���<9�	T��*��r|
�7�.!IG۠	���1�K���猹p� �B���20˸#�u�܊��g�� >Y�
c��(�a�'�4:/��5������_#�бW'@��
�d��m�=�T[����McMgp#ڞeN����".&��M�Sy�I���-�̐���R�05'~2�hZ�{w�Y��,{�WI�B��h�2E��
Z4!����8����2M0�����/>�����rHf��k͐w�֜nU�D�
!���E��Lk� ����?��̨Q��H<;天�a�  ( L3���n'[�w����a<�C��d����E���X�y�Ri��>M[��l�`8�/�$a��jn�Wv��>�i^J���$:4K��I�Yk-��C�"q���?�
��}e���m^+��3�F �������,ʂl!_�<|��uT�����(��w	�u��6z�ݗʌ����Or��|h�3΋[�BG��|������������D�}��b���&�e��!MѲJBU���{ҋ�*�1�94����y�|R�����ѕ����u`��q��;�s0$l����4ƀ#w n�.����_�N@:&����r|�Z-��o���׮��X̢HH�!B�,���+��W�f��ѐ�3{.�k�qf�J=�E"�۞u�	���ҕ�i�N� �Q��΋��֑DJNK&!�ך�����
�j��Ÿ�T'ɩ8;�ȥ�����'�̬�<a��z��L��q72�(��,��ӓ.׼�vFO���m�u�@��a�:q�� L�J�yt�^y�ڠA�� =�2�� �$z��~��[|lE(F�p�@af�Ɛ���+�C�]���-��R&x�I+x�B��s�?V��A��>�_��:�I�s�1������I�e9F����NG�M�0��J(r�a�d��r��\���#A(�j �Q��V"VW�[�T�^�	���p�o�O�s�J^t� ��$��bu�2^���'?n/[L�T5�)/��G�c����`J���=�D�/���؜�UO�+�~���~��
n���MA�  ��\�g[�:�> 4r�:L.\?�كWq�`��RF[ɔWՕt9����i���	5�+�3�����|�##- /��j��J���s'�yq(�,�d�3j.�M�3J��r->����5�j��Sʸ�˨m5�VdPBO��3��Ft�J�dO�N=�C�2���ӥ�wV�zJ�!>`+@xJF�e�A�� ]�!Z���%4�'����z+� �� %���ƋE�	�h����}�w�4Ƭ����B	�����ܼAL����4�t@��-�m�.�����zm~ǳ�3|,��Fq�?���zȮ����
Y�˻oy�bA\��J�ǯ|�����T!�� �оKA�I�ct
��ԩ��4�ئu�?��g,3Oiw?mo�:}����#[!�)�d�j*7�Ϳ��Ehߟ�ǣP�FҘ?�Y��bS�C�`���:�P�BƖNf2�U�v��p�6
2��K� ?ĸ�v�$���-J�Ě5b���I�T'�,�����<��:d剘y@=�E��eE<%�;D���ƁXTH�F���\��O+M�1� :�+Y`aOɘ��<F �tr����_���m���zK�t3������&�e['A̯D�ko������NT�$�R�]=�'�@��)CDFЬ}����=�b��'��6�Hoi�F�\} �v_��K7c7i4�4�!�G���3����U4M|�j=���:������.�݄l�9�ᵺ��������/��W�e-[DF�vy�7У��D�\����o6wx��s�$���~��"P���dSm��F�O��{��ҥ�l+�
�ܤ��d�}]�dwn^������f�W���a��Y�2�˰T����=h{� Q�)<΀.� ��F8�}ߖ�Ŀ#�r8�l���H�0��A��� ��(�T�����(^��+2�
��1��=��A���MЍ�7�8�҂
�]�~Ju��)�߳�A:��ңP�*��1�>�j��D}��ɏ������d�uOV2O�i�$\�-W�Wy���>�������"�D�	�Ȯ���ŕ�__9��k@�߀�)\0n�Z$X�&�0���k�j�|�1m�zaX3����6�P���m�Hܭ�~&���n�╘X�p�:ܪ���kH丠]E�e�� U�oNy'����gF+ad&�L���{T{�c��;�'��'`��97r�/*TS��J:��S�#��Ǩ��.���J���Eb�IV�fX�ҥ�tA��?M�����A��NV%~��y>�sW�G.�j��B��Gm��^h"J���j�b]�vf�\�����ɡ	���L?��`�@Y�3�f��������9"��1O'eG�t�mI��8M��3KȬ�������*�w��QJ���"4Lq�V���^�X�{*v6�p��L�t��J�v��1�^H�3���� ��� �o���(�^їWT�D�{v�Z�=I��4�T��)�d�>�c�z�L-D~4�[}���rFg��ZH3��`R�S1yUKZ�O�E��A�������H���*ےP�N�����
ӡȻ�ђ@Z9����K߈��_�K�Zq���Y���ǰL^xA$3ig�谥Q���k�y�L��"�`���.�`���7�"f��`�AI�p���b2�j���k):�z��ݍl�c����r�� �S�"�'/��N$����OgL}�A ,8�ϬiC��85A�*l������>j��R֭_�H&�m s��H.�T�3�t�w�D�{�AR�2h�e��/z�#��,r��H�T)@#y�Usد�sf'0R8���q����Q��S�XW-�	N85-,1Æ��X.��4!VC��@��_#���.���ۧ����ghSĝ�j=���,}��:v%���k���ǹ���oVG�x��d��;e⊺=�Q�L��7:;���cp�tp�;�K���5G�5A:�B��!�?������/��-������(~�7��CA TB�m��`�����
�԰�k�sJ�yke�$�M*qrTº�M�*Ѱ(�9#�s��h�x���W9��e�
��ڸ�ݭ~ŧ���\�KK�p\�R&�b��gI��F��7?�`C�Jt�����M �͙ ���OX4c�OU� 	|p���lo�1�l�|�>tH�Υ�X�.�O/[Z�Z�����~��g:�A���m9	��f�	��x�����-u9�f�B���,����_B�sV�W���®���	/\n�S������T$9���}[��)���5p�F��~v��*����y�tű��A�[���I�'�Hk������8"�з����-� 眫�*��[��Փ��W �l"0��g�=��\�#����W�,�ֳ�& �d����E��c͏Zq��3ָ4x�E,hJ�� @�""C�Ū�cr����`���;�T�[(�_Ip$r>u�ZX*E�̜|7�'���\��N`��CKn��S���@�MH��І�^D[a�]2����p��D��ޚ
s��>���Z��h��Y"x�t�c����4�8�6��Sx8Aɰ�.�>/�s[*F������F�ۧ:�z���<Ӭ6W)�H�J' VR���b�nI�;8Dq��p*0J�{���U�ۤp*
r�#����B�;!��E�~����O�m�Ż��s��Zy\�=�?a������^�A|GK����w��&p��p�=�,=�pﲘ��儓������8>l%cE0o
�×iK\�_�B��3B>�ɷX�U�~�����O�F�<1kz�x>m��������/bO��|!��;��k(�+#&U��A(��ȡ�a���ы!NՁ�[5G3曑��ع���K�c�)�]qK����:�I�BO����b'q1CI�7noza6���׍;{�}y�3��頻�J�n�1@.c��ba`f��[rK݇[f��	;Ĭ>bo��"n���0	bL�����-j�"��T,��m��~�\���,�\	(4��]���U�������D��F�����o�	����^ņŌv4MO[��q��MX�?�Am2\�w��Y@6yք�,����E��=nq@8|j�9�u�@�
��.쉕�A�	70�'����VfcYBu1�yeOZQa|&��42M�,�&ݡ�KVD�f�4��v!���֪:�͋��+�2Rk�,���~���I`�`������Do�_�W�C�7���Ά�&X�F�\E�����P���vB��ĕܦ�,�R�������x0r�(()��08*c���Q��,e�Ә��;ل���m�O�E��qJSKqZ)W��?�A>��Ϋq �Vc�1���j_���CL�?�PL�R̃�c�8�Dc�9W� �I� �Nqy��I�el͚K0GU�n��!/����^��a?\�b(��ʙ�	 �Q��?�-��4��т"��S:�<C�#�h�x�"�����o�ٌ�I��x0�x��C'��7v�I<+tlvU��-��vQφ������6t�W*JP\[5y���^����|�q_�Q�
{=�4Lmį�U�3|e�9��62�S�(�DۆN����ިw�SmL�r�����Yr$�Q+5�wӃ���K�1�N'�����(S�U��s� �2K��Y��in��fW��r�}9p�W˾Hҹ�̺�&�,/^�k1�����,���������s���ev� bbeq
W��1��>J�XN��:��!�a,䧝�ݿ
���V���8݀2��=��Q�q^e�
A>�E´7�La����N��jp
g������.�v�f.�6�<8G�T�m�A�8O��8n����G���QI�����2���?���}-,��R���;"J��"�x+>�m�Y���B\WG[|T�3�m�r2)b�v#�7m�Pnt�~a�6'�#��[�p��Gj����}��*���r˾A=z";j'�쏯���|m�ҭ�a/����۸o?��춶�g� � >�XM�������$�T!�/��Ȧ�4�TLXW�xL�2y��R\�׫�����l�.
z��k���������&f�#�ڛ�de��9�U�s��e�}3����u�Ўq�c�JC����&�]�c?pn�plz(-�dFQ�^� ����zn�"y�c���H�}"!>�~���9
�W�N�Vk3`G��Ľ��ܙSb�s�_������(W�r1�����A�Aɕ�d�ķ:7��K��+��7��AL��X�(�V
�[D��	ɓ<������W���#_Ŭ�*�c~���"�5�|
_�E^`M&p'GQJ�=���\�ʿ�D��m�u+Ȫ�"!������"��ug���%��kE� ��T,�C���:) ���'�ɏo�V��ƨ���TW!�q���-���JPHʤ�ЍA�;P���}�4�j*�����j�����u�z�Xw	�y���i�I��fn7wr�e)��TUU�za1?<_���į"B��Gꇐ7|U�>� %�V���c�ax�ߙX�b�A�q>RM�"�2̵��$10Wm�����`��K�\F��@@���}�h�W�^}�:d�I�����WA	���@1�=;c��0������ >
��|���Ő�7�@��U`\5�g�Szx6J�TjF#F��k��^ɛ�[~���BUq�7�W�i�q��١�ޔ�?�ÞR�
����3V�ˋ�hN˭K�뛨-��EG��W�B	����A��0�1%��dΨ�~3;1�_� �x;���J�-T#Vr�JE��B 9���֠C&��vc�9����B�o	
�����]D�>vb�E�LNN,��8�w��Z���^�]��i:t�3z�jOد��'C@ >�(��"��ƨf��8������;>9��1O��]�c��?�=�K {%Ehc2��j��]���Kkd�ef_�,{��KPx�p�tx����b���V\5]���^R���[���"OE1�����XV�[|�|���Y��Ѫ��YG�\��S~d�3��;�F�&��g��7�7]a�z3��|ȉ77��XsYQ+�dX�ɹ������ޯ�+�צ�n`�p!��TMB:��fЈ�k F$%^@�%v B�G�?�A�v��"���(��N=]�U3fC�l%��!���m��[+#�?Ϭ�i�a��F�p-������Պ>@�~<�(z��+���ęJz���Z�]Hm)���X�ܔd���{��c��3������3�7|+6_RW�E%E�v��ɾ&�*0T��y=Z߀��ɀ�v|駡F}h��H�7���Y���3'lێȧ����v�S�	3_�O^���d[�B~�����:�Y�Nʖ���s|c���C�� �L�8�8j��fs���)�P�y%IGI�!�}?�I4���*��EA�^0~��/�����(� #���8Ygy~F�O�Zۛ�?q��z�k��s�	[��*"ؤ��I��7�$uG��wI|���[{�m�����K���#FH��	f�n��`W4A��{��XO�¾��կkٛ�� ����1>�����O>O�̇i,3��V=%�����db�� P���CSc�k��@S��������wX��,��i��&v��.�����蹛:���)V�����v*Ζ
�mibf�7B�Im@ڪm!���l�=ߛ��,���~.��P1[��^[��:��B�O�ZM�&��� WG�X!���I�:0i�R�L��cH�C����i[N���aF"�xě�W�TB�~��AnI�N�S���z7J��V���ۑ<%����=)ʬ2P�[Կ���5�40��d���dHIՁ-�VϼJ��x��n�h#����]�A�MG]��Oր`J�����0�f=4l��'%�� �$Klb�h�y���-�4+ �_Q�`2�	n��q&�d�[�R]5"�6��(\�T�%ö�d�E0�cy�F僤p]� �$y�h��p�yz� N؁a2�QKI�ߢ��ش���zO��}�0Q�#�p���=-ߏ�Cʱ�_�3I/F�~������Ƴ >�����4��K��`�W�*>1�5�(8|��vbῪƴ���f��$��nˏ�~£�J��N�u�>a�@��v�z+��z�D�.)��~!	#!��_W��p�P�����%�cJ��B���x���w�:e�]*���7�Κk���4-�'$��Y��� ��n��E� R�^>���6����擯n�ǨNg7�E�\�a�_Vy�a�� �+ �&��J�:���!�rW1[����"����]&\#���Z�l���JHX�X����]� V�3Kխ�8��Ojս�ʏPL1�f_P�G{b��a"b��I!~�s�W*����e��F�36�K[ݬ���W��j��8_a����8v�7{=�/��w�i��֛m��Y/"�g�ǡbrS�I}3�`�Ƿ"��e��EF�x���`����'.�pv���N�s(�!>5�GO�ˣ�5I�?v7<UO|Uu�dG@���<0�+�:8ݜ*