XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f��Ơ�!�6,Jt�͡"��Z�`�3�|�d	+?g��@��u��#܌���o.�o���Y�Ii�$k������z���|���F��LX�!iU�^�'-޺/�ۆI�M
OXE7�����jb^��22fI4��Ni�*���s"_HS��x��,
�d��a��%�	�7�O�:����i/1Hո��x�h]^���J��2��d��^�f�k��ަnC��Y����H�+2�6̀���N,(��*��wn��ՖAѽ��xݻȌ����J;�#����k3������Ӕ5S�R���-��X�Y}���P��fR�T#��OeO9������^��x�'��]B�	�� {9Ȥ�C�ѝ�bX�Ӏ����|��^+ϸ|��m��1���P�����I���&p�*��x��w_����$m@�|l�z��m�	��`A��"N�
��s�5w������N�Z3�Hr�-�B��a������Fқ]=d�~*�C;�{P)j��ȡ���:����1�m}#�Ĥ�Ԭ�
zk B�%ѫ�����`���ߘx��$ꚰ���`����_���=�:�Y�V4s����"����r)Vh6�H�͊+H��&D�Kj�БH�y��y,�>&�f��EB���Ͷw�@�B,$��4k�6�$���aI�9�����|iYK�E1۬1�%�r�m�NΎD�w*?4�Yb�4�}=c�dJs���{��vc���n���,g�oXlxVHYEB    291c     cc01�vh�-���Zo��%UZ0�nڽ��_�P���^n��3��������F��9�NGF}s��6ҟ����0Y��y���,�e`���u=5�K�'�^@K��|�%�f���.�G>�ʝG��y��M_f6����x�����H����U>���y�3ZY*��K�)GX��-��M_Y��-��H{C�1h~�-J�л� ��}E5�s�SH$+��,���|�C?+��<�#��3_!��Epo�+e�3X��1ӥMS�6��������$�_0����j
k	��c���<��ٗ��������9��'ͭ���Ġ��?�L�jjE=T�.}7+?���v¡��%Pײ��r�t�����������>��Z�Fr�4�@�����pCIB�告3�/�q���ItEl�w� ��)TҶd�7�DZ�ɥ���҃��C��|lƛo�Z�i�6�'�y�)<�n�~�D��u���6�gѣ��	�K��(b?� ���ΟiY%��?y�c����`[���nI����hAw5З[@;��co%�=&0���*��uϚ����	A�H;|���=�}`tP���-�p�%�{�F�;G��G�te�R�r
�1vMj�r^H��_^>	/���T�z1:�u$���6=E�ky�A��X��"q1CY�,�Z�# �L��^��+%x��'%�:4�e6��ī�.�4^U1<��J��*� `��.����s3@?(�x���>�$wɂR��Uo�v8|k�X��t���FxW���Ul)n�#����dY��ޅ��>$��2��?8��J$L
�z��\S�e�b�H>��"H��P��=V���m6���F�Ĳ�_�|]G'%���=�!��w��S���,Mk=sF�@�����x����z89xB�`�7��u�#��U<�����d���O��,{����~7x�I5���bͰ�w?�_+�˝��}��V۲SӶ>���u8s���^c���/kDX�շ����D�1
9����	*��|�yv�����(��g��E�إ|1�/t	��M䆎�&Bc��K"T���q��ƍ�U�M��:v�,�)o&u������w~�n��:gT�8M@}��a�g�������+�z"����o�zKh�
?[�[)�Cn?����`�='��&�b,JZ̵tw~�(yP���҃��i�*Ww���Pj�SS��k` ��:!㚜��4�Ҵ.U��`���g�*g�qT��΢ ,/�?_z_dc����qh�7J��:I�9J�+�.�<�ބF��=3y����)��Y#'�s��'i���)$z=7K6�4�?�{�?fmv�j:��{[��%�/@P��a�<��V��/��/���)X(ƛ��������`q�R���Y&�j�Kk	E"���F�98+*6������{���u���O`W�yh?��.ʸЙ+�c�
D�j �i�$��I����y$k-x�;�2>D�H$u�D&��'"�z�2 &�Px
s�`�ٷt��:i��)(��;
=i��ksXl8]q����J_&*��Z��j��܀\(�+X
�����>�9�+!�%J�g��a��5JGg�;'�a���M(�_ӭ9d
���b�����"F?j���D�n������f�n*`6W�41�KCXhB��F��@�`�do�N��*�M:Ε��g��TӸ�x��q;�G#_6�����+�'{kN]�j��]?�ȜXȄ�Q��j/͸���s���҃�G1��>���cMI��6���W t��F�3����C^�q�!�E�]�q�����j��E1���Ia���k����EvdX!o��Į)��Б,堁��M�n��VF��p��̘��&>�>""@��O�j���]_�M���V߷%��4�M}o��Цt���#�n�B��r�P�P��=Z���&n�����n�J6�v���N(��"�*�[����
|�yM��_{B"��z~�|�n�� l!��ZS�o�c���/X҉9e�l�t����0o��ߖ��ȋ����m{]4�y�v���
m3���=7B�����su�}����2��Bc����Vo�f���;�D��E2~?��KV��RK���rJ��K=���<,�^r�Q��ʥ�2� ��l�*ն�5�����湗U��p\��pQ��n뫰��B[�Af�� �0�ﵒ����L��!&�U-mrݔ��b�%M��rOr�)���^[��Bmďwh�w�v�,K���|���J����.wKQo�_Y|�/��p�<L�d�0�p=�JK���ٯs�|K��1�(U��f�zj���6��4��Z*m�v�H����� _D�+u� ��$��0�%�O���R<-!���}$��{�oN�Bni��R��r�Z��4�u��	_���[�X���M�;f�8���&������ʽm�P���`@�բ�x��+�t��n̓��v�Qr�����s@?�q�N6��8G���G�[�j&%��W��Z�K��� ܗť��R��GZ�����AЗ�������m�
��w��5V����~9)���#�	*!�Q��x3�/گAe�W�c}<��m�X�x���|��]��b�2�Eu=T9�@�FE��͡�]�$���=����fPĿ���<l�F��?@վeΤ�y�TM䜓׫�
����lȵ\ˑ":�`+�]��hSG��_�6�o��ߑ�%́�y��Tp�Rm&���7v�$�$z������$m"�㎽o�ÿ
�<<��2�׃u"������ߧE.v��Q���,#�u� ��6��7��yk:��ϖ�o�7֔=Tf���j�ѐY����M8Y�V����CC9��WWZ-&�G�Su��R����nz>c��4p�ĕ0��Y�/�h<�6�f�V�Ao��n���,?�/׸�ŧ�K�]�Kd9���E�e�2�Ut���5�&*@O�4�6膺A�2{^ �
�?~�f�]U�m��||ft�v?]��Tr�ީ��PF���z�,��}���X�\E��
5�Z�gCJX�~�d�����,�I��z�l����@�cߋ1u1E3�C�Euh4�J��+C���F���T�܏hϣ���>��mŏ%p��j��[�p��l�s���P�hXh]�FY6/��j�b�� �~��/�7X��^T|��.�!�0�i��N��K�>��m�|� LWzJ��+/