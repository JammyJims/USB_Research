XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N��\=�B�D��z�;X�I��ɷ&�m�݀]�8պ���$��^�o��֜�n�#K�f�XM�m�zߔJ�Y���?�)q��r��`|�g�G���.�<(g�,�k���.0q�dk�!��"˗6e�[
�������\Q�!p�z&�^��A�F��k��NU8�ʒ���|��3I���"/g�j�yԍTf��4������$��wTU��Ͼ�kf8���\�L¼�F���@�.I�Y�g�������3�g����u¬rU_{�yh/<TAe]��b�9�ɇ�G-��Tg�\c`�{��}��/���9E�⡯#�c���d
0�ERF0x�h�˖�Z����>���iS�U���̀������v���W��!�,�����[i��ܞ\�����hN�XU��4�i�.�ed�T7�4(���%Q�qk���A�{=�pc�b�%��s1��5��]S6�Y���u�{~�J�����#���O����ic �^�R܆���T��b��=�]�����I�W\&��|�Ρ�]qCo悿Ю���5�����.mXz�bK�BaY��t)�� ��b�ȕ��*2�o�`I%y��>*<y?�R�ԓ�%�k>v�O�v��ነgW��An��2S(����|�����U�UՓmj�Z�����H�$�����v�N�	��v��.��0���S��V^F� g鲓�H�N��T�r�XH�fT_ڀ�P�p�V7�xD�do1��6HU��{^-�~������\��=��Po�XlxVHYEB    3c4c     e90ݥ���8���I�	Y���?*b�-��K!��D�r��>}'CP�!!����u�t����_ϒ8��=��9%mU��?s����(�ƃ��X�����(%6��b0(u�~vwSx�1�ѥh��ȯ��0�eP��]���mR8O1�a��L��;�jdV��PY�!R�/5&9�w�B��X�c�NB����S�9F�,�y�e-`7�>k�����b��t�V���H��|D��������c.��;h����莳�٫�`7 I��,�C�׾�O����C��\�0��{36P ��5n';I,�oޚ�1x��E��[�=g�^�{�1q����E�r�TQ��߄6�&�d쑊~��~���~'*[qfT�Z���ҰӬT�h2��.d-��DW��<��\Iݣ���l�:,����r����:Q�(@�^�͓)��מ��M��O�2��9��������W�!.�C�|�	��B�3�}�dޢ�'��� �[}�hrdj"��C�s�M��>6n?�Z����+�r���)p��9T5��"�9��Ғ�j�ĳl��I.o��5E�������e��`�S�#�Z\ ��Q;�T|�
I�и⭟v�� ����/,� 8^+4�E�~Uզ�q"�?�Ag��0�g�Ǭ�<��G/��5�ͬq�u��v��'u� UYA~J,�D�]]����k���@X����`H����Э���I���������ݭ�mQ<EQ����H�ӸD3ǂ������yF�W/J(E��¾��fJ����H�MDq��ة����f�$�'��MEco��+gB�[k�~6�N!R$g	ѸfQ�4@���Hr�,�X�T=�O`x�0B�r�%��o�Q������-��
�� � �*���KJY�C�=kv��ǣ=�?�K]s=}S�^#!�ܪ0��b;dM2��&f;�|E���J�#�'Y���`�eH�S.���(§��p�~��}a���OTY��Y ,3�n�X������a��'����֠�	K8W*�^���x4P���T��C��琛�=g:Y$'���;�(�v���a��`����<3�՘��{,+C��Y�&��V�D�K��R�^v��Z�ݳ�^���/�c�A��Ēl�\�&迊C�u=%y�I�x'L�|��Qi��tH�c�)�Q�NR�p��5\N~�XQ n�%0?!��t����R��� {/��pIxV��iD�p�1k&5�qY�ࠞ�:�]?�F���H�v���\��˖(�y�x�3ˎ���
�}`�׋�[jvn��]��b<(��G~�����v���#��`�����ڶ��.hS +�W;x2���O����n�֚�����w���btt4:�i�{Ѥ��|����9֜�2��`�P��j�PXD���ˌ�e���j�,M}��0��ZR�?�g�+�<���W[:�.�W������F����	��E��le��;�k=�\e�4�0�U�DD7
(����y{3��绐ӻ�4-Y~N�Kz`�mS4,O_s���O�%=� D`2�"�
�ܲ�7���*��Ќ��0�grd���i���*/鮢���6Ҵ��a���Ѽ�hLo1�Z/s2bh�O��ҕM�5ɑh�A�2)����������NTE]2KC�2u��P)�Ј|�&,Y�Le��<���ⱜ��=�G�=%�䣮�1d|�e���?[�� ���6��̚��P���T"Ǩ�yؔ��n��4WW_b���_/��� �	W*���.;]z�����'��;7������z��%�Ӽi��O�;~�'{��4�7�A��l���$���+������_>�E��!ٛ��C�W��r"�y�)1 �[�����ҥ�i܏��RfS�����l�&��������ϒ�l�U���0���)\���\SD�;�[�g�����)(q�۩����G#�����6�]ܪT˹r�5��ɣ�~�Kk<�\H����%SK#S�+VYE��^��<K�oÿ5y�h��O�0�g��Q�R�:Z�e���3^a�,"�g��UF����Z6�����������6qr37�;޲*!��$/D1ey0�4�6����$1�M�j�T'kN�����eO��	�z�
����+����:R����<����4�tqg�t�ذ��6x0�����8qf�	&8=R���W��:�^krH���wRP�6]s!�Kz>߫A�Ƒ��t)��5Ϣ�??i�'LG���H��l�S�v�8�%D���c��Gi�tpo���a�e�y��Ȝ8ݞ3��>rm�F��Dq�>�0:����s��e�ȹZ��
l�S'�D���|*�V_֚'�:�񚀞���:�mƇ]��F;�e�������wD����d�t*�B��i��b�_��Z��<�͇q�M8����Ng_�����7�nx�G-f\�^��ɜX�̀ѵ��c�]��Uv��n�q#ݱ>�BnS!����u�l�?��:��\i%e�zFR+/�WK�c����%�c8�B����O�_��f��-P��Y;	�agE�ܼ(}� ���BM�Yj�{�C u0ΘzM�t ��[;Sh�@��.��	�2�^�ڪ���������"_y1h5�:��?;r������*�.���=�{�-]6*r���� �'e��S�D2LKZ4�)pۊ�Ą�M	K�dB�;�FLoD�b/�OK��e\�ע�A��:?i!�e�~[ObLj��(�7��Z����1�I7�W"�,�NEa�U��a�|�d;�J,Eb���<.�rˏU ��Dj�'GCd��������(cU/��f��[�3>�H)�G�p��s���j����3�3�&G¦c�
�J��a��5�3�l1�?t�;C�&�(t��ҍ����LT?Wy�GR���0�?�7(j�]����V5z�Es/4g��2��â.(,��29;��u(�P�݉�eDy��Gvo��z�*!Ш(�6l�AЈa06��]�?&��*|�$��&:r d���|�W�x3���m��6�Ć�ɗš^ѩ�<Z�P\{F�催r҈)������XE�ƖhB��@�����ˉ����Տ�ï�����8,m%G�4�
��\�F �c2*)�@����T�aax����r�4ϕ��@+S0�nf�������^�\y&�%n���_�<*�˿�X$�mt�ه��<�x:\�Xp{����t;�o|���]�<kZ���)���J�4c�vҠD�k>���Ʊ���춴R͋ųFo/��������3ծ;kgmG�֨ A?�&���܍�iܜ{x�aM�d��:�w���1C�JX��7)��_��������e��q�a��=j`um	Z!�>��N����Bg|���aFI"�!�j���s�h�?(��=-)�M��Л�"��R��.��Da���F�o��� �IՒ�:��՘,z+]w�]밬w��H��r�+"u��/v��2�� �U^��o�t����C#��������N���}#�����[��r�� �Э�o��\��Z<v�X���ق����տ�V��Y*7�V�K0���x��(S���^3�\��o�$W��\;4���[�Re� �'�D��G�M��C 'D�Tf��17?8�V'h�v�J����d�S��