XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��rx+U�0�}����T��H�o�8�*�g<�v,���+�fD�if�On�P�9����w�r��_������/jx#V\���)��C@NZ�����uQߦ"�6�}���6;m���ǳ��.ӳ.�2�ˏ��x�; ��mW�]�!�~Me9cF�ݬ���L^��H2_��;����i�h]V�Tx�����Ң�Z1��$'4'|����`A�j�ԯ����=G�tt�P��+}ˑ*���(���d��܄�}+� �d��O�ͮB>@� ��N�^�BT���,�� �Hpz�T~ֳz4WN�Ģ#���T��]]}�=�N�{�A��q���nʁ�g�.!y��P&�R���\䢫�M��F��Ѹq�m�P�)<I]q-��C��g6��o��O\���yJ� ��\Ե�iߥD��a+�u�p�,m���C#�m�X�ьU���~��}dQM|?.;�&����B$L�2��*��M��0�ÿ�
���:5��I˧��upc�:��Y�-*v���H��� {�?��Ey���9�a�eͻ'��l�mca�e���.q���hֿ�yG�Xx
�����:�uV���ڜ]��=�޲4?�r������@����Y�� W�����.�@3��m�#���,HPT,)}^�<�ya8~��K'� �L�{�Ò��~.]%�����V0�>�D)�����}J�a�'����-�U�d��n�FW1�:q���J��g�<�|�Ϗ���D�\#I��C�g��XlxVHYEB    fa00    2e20o�;��Jo��֐;X��sl�F�,�=�N��!�w�����v3i�B��D�)��*w�	�0�"9�a�{b,?y�}ѣۣ|ɹ0�kL��O�T�%�ùKו��W��n���E��e�S̗d�9�ľ����*G�?��_���5�0��Y/�ҵ
}��8�����u��)�!A�^�|��g�v7��ǎO�o��>��ȯ��2�w��}��iv��7{T{���̕T��E����(�H�GC6��Q僂�����쥫�5�Ft��!LL �k"��(sv�	�{j���Y�*��V<�WFH%i��f�{��S�>S\!1�@B:w1͒���=4Oy�)K��M��|�6{�T�1������bTu�u̶�?@Ĺf}�$z�0���ݢ�#Y
'jF�������~�6�������d~,�W
������f�H9�,�ؑ�i��2�cMע���r[qnb�0�F2r>�,y5��A�1�^�^� |����y��v!�W^�p�iW�*r�mvߒ]�}
��C%��V���@Ѿ�� E�-��K�Ύ�.�\b#Ns�C��F����V�о��yZ�����t��U��hx�#��� Z>.��8yP�pxm����,����P!?�P_�V�t���9���]'�f��9�+\�gA^��T:��S��8J]8���qz}�cvfG�ay�RNԺ��k�+�:[c��a��������z�^�� gw�Rv���6�H��9���Z�c-������Yo|���j�(n�}�4�A�ƒoU��㞑����Yto��]��ZU,�T����r���H:wcT��C�=��+^%���qG��č9A�
�nY�wD�Ρ�� ��7����k�V7�<�K�.����:�9\��;)a�#l{Z�J�<����moH�Y]��
LJ���5��O�톾&Q%�B�0A��!]T���M�qg@m�	���H�$Kz�``���<`Z��/���D��#�ե�{�|�T���U�S�d���^A����j6Q��9�����^4���v���M�c0�w
�:�M�47��\Tݽa;��}���"��nݨp�ਟu��$���yH6�$��)ҿ� ��7���������d��_ur��(Vs���0Գ�\�c�&ݧ��d���E
�����A�5������ }�~y�a�v4�&�����ʯ��\ΐ#��?�W��ch4n�Ū�r�҆��:�l���:!42��4�*[�?���o��B����x���o���f��,��~�i�ȸ$�a��_(	�ћ`C���pdˀ�g�ۤ�;���w#Y6��d������V]J<f�6�
�����������Gz����q�Þ �4¬�ܷq]�E�J�8K��ⴅt$�0	
�X��*��3�ufs�vC��m��6Y8��VՅ$�Ϟ�#M�2��ژ�<���[;֧�Q���V��)����cZ~��Ln�ϥ�i˳���ԧ3a/a���ŋ�1xU<����0��O�w���!�J�D��(u��3���rC��J0d�|�<���Og�놢�(�A������P��K�FK
"J2����1�[?��dF�CER���4,o�I �����h�pPъ}xU)8|�q�:}�+�P���v�T�0���b����cY�Z�@�����������9�G� p|�ށ?zN������a�H��j��ud����_���/��-,��I�@����� ў�����Z��=�/���rW����"A�'�C[C�8hS��˝V�ذ��?�Sҧ]��!ߗ��� T�z���Ы��Df�EP6u��p�-�l�9�_f9�Χ?ոS��yi���.d~��p����PDv
����JZ[�2s��~`��	�2N!����ɱ�G����U��O4����8ޞ�U{CƠ��T�-j����l�oW,cD��=�U}_/��P�U ���Sk��U#�e��HTȭ��!�"ӈ
T��ݨ���������? b�H�7n�`��Ơ\�f���W�4������)`�,��>@��k"ؙ��g"����{Ў��t?/Q1+;�����vh�ȡ�G�㜓��%�~#	Y
�C��o	_�o��E�83�R�]�\�����t�'$�\���
Cȋ�a��E�M"ʜ����4SŨ�]�WR����p��~�!�U����f�VTI!��b��P��2ГDj�=1�O�Zv������AI?�]G:G۪m&F�is5��L�fu�JZ��]�ρf��AL?��ǂ����Al���4���|��Ά�-�!2֯�C4�
gRr���5>&�)|�|�3�ᡑ����R�ibK!?������o�2z�����u
!K����YD��?�eK@O��<�'�4�!j-ѥ���V�mp���T>R�-��-���\�"07c�a<�t���k��ê�}O���K	I̎�V��sգ�]�1���������>=�_e�uA�[���tY0G=N�ǉ��`D�7�sB��s	=p��ҭ?pwB 7�[7�gf�[��Cϋk��K�'�k�n�a����2�S�C��3��d�OrK[d��
9�)]�,
��0��  w�m�$1��sA�	�@��z����!.�Ms����vM�:�Q�w�w(��s���a��^q/��/_
_g�!�c���ѫ�i-�qR�4v�m�|��k��#�D�鐠�����T�UO6P� R�����9e�lb�fM���y� mO4>� �r�4�=��-�ג� ��U;�7�}���}b�f�Î|;����Y������]r�fx"�bj_�̒�mM|J+U�f�Ѭ"�D�j_���Ke9�{���
>ӥAv��9g�ȔK�Z��;SDp��,H���@'Jh�33W� ��
'(�y�2��i-�i��I��`wZ�$�̓�o�����q��_��QS	,Lk&�-m �/���>ur1ۋ֥\��O{�D;R�<ɝ)\��ĺ~�y<��K%��kV�[�J6�O_�r���[�x��H|��w�)^�,Ǭ�ɒ+�[~���s��ǜ�<ΣA��iX��Gr3"Ty��3��An� ��kY�=J�8y^YE���1`T�Z����b,�ge���ZČ����������OYu��\%�%bk�9
�Z�ݛ ���X���l_������F�v�G�����]H���ڛq�����C4�Rb��j�S��4�{����-00�*n�|Ϥ�O�F�cj�Rr޶�g%�|��K���El�0.�wFu&����7�B�z���X��	����K�[���������$����=i����5�?���EV�]��r�u<��8l�<l��s�3��{yMӐ��j�0�'�9 �t{
*x���Yu�f�W�̞��D�?����r�����r?�X�ϑ���E����z�b����?�������el�tx�?��=a�������J�m��XN_�P�JK��E�q�V�}�� �2����B&�Q�߿&3���F�4Y���x���T�����;��ѿv��P�(���bް-������e>_λ�D_`#L�m���B�h�P�r��Ò�e��l!LR�ݽ�?O�S�2���zC����m��ZZ��!��U�ȿm��È���Z� �%����h����m)iYۺ�1-$/��t��ؙ0)\`Z�$!-#�U�ެƣXV	X�Q���8;&wL�[�0�����Z��+3�2I4��J¼�Zǘ����Xz����{9���h�=���L'X�}��UO�<ed�_��xz�G�����m0�(�e�6����y~�م�J��K�3��8�غI$:���*�{�4ME���d�	�z!�|��4�W;��mףc-���}Ďe�Pj��)w�鏞$&��μ_�7}ּG>��|�~K�Hoy���JOG~���U?���TϼA��.���i��d�fs�>b�f�FY9���X��2B�x�t�ݎv�)���L=�`�0S���}�,r��! �q1TF��i�=����O<�]u0�'�2s���v�ZRU
�2k�`�]�7t���'��~Ӹ?�*��^Ҟ�߭���K���Sl��l�-*e��lS�pR���Y����`�0�Z}d%܆��0F�d����ē����c�x|
�4����o&1��t���a��g�Hg_Z�]�\x"А��Cf����z�=�.�Np3����3zThk���>�$�����-����y*ox�"As��o���k[)�)v�2K[C�}�Z��)K?"�����dɨ��m;#�����&Ԫ��(��ISf��4F���b��ca!����Ȑo����KN4�~U�7:��k5(ջ�ڀ[	0ƅ�nJ34�ύ(.C v�!CAҐ �'-dQ����͠;+����(�����୎5�48Ӎ'a �>,�%�)�따��J{�6�C��VK��������
�I.���}_���t�[�X�F�\�;VP��ۆ��+����1�r����$��������AL�6���7���1�=����{��FK��T��e���P���D�Զ���^&�pn#vfy�9I<kjdy���,To<#��k�`@O��:2.Dm�9M G�0W���7��Ɯh(s˯�K�0#H{}�6�c� ���9P~ф_��P�l]�ᔴrb|��V����p�h��Ea�`|dD�[��F��d���|�.�W@6WN�ٷ���R{��1*,��@��jI1�n���[9y���j��:�ͯq�@������!,�_R���.����Fs�@;zwb��"���RQ�h.���Ӣ�V�K7������b�7�&�`�P!�xh-�e�p���K{{q~!��0r.�����
γ��c�^Ǜ+�K۴�Ȕ�B�.�����6tx�=,�����E�)6�n' b�4�GI:�f)+6�g�=ڽ��ѓ�w#�����@��}qg@�+0����Չ2�t��xke�5����{��:��0%8Fb��7h�O���j����X�  �^�~ض��-}�{d�� ,���/���A����ԡ%���)��I�2\����LJ�(����#�71vv��q|[V8�:B�n����>�b|���7����+y�kr���z�s�����MpՓY�s�F��nW6{1��J��Wb�J���NM���82�E�$��u(*ޥ���Bd�h���j>c@�{����<_������]6���nb��ltM���zO�����q̿��\c0���UH}��Jr�,�Pv6Xzp�R`Uw~HYė�c-p =P�Z쑑o����V� ӛ��m��ނE/S���x��sK�Vr%�Q��'�o�\���'\���+�c�
��*ѹMc�+@��Q
F�xrԞ�ƿbt93dw\i��ԞJ�f�#� �5�̖C,��{�`!���|~����,2t0�<�<��W`��oc��'�ՠ�� 0e�_����ǯx�gpV�d?�<��n�y�iTXӱ����������Ä�̖5}���ǣ�f�MCQ�z��Q9��O���o��{���i��(5��J���Ub��Ƌ�ig����[�=��sWu;�ZJ��x!J�%M�}�^1���Iw�v
��<�!���N{�.����rt��yR��u�d��������$���!5{_�A���BL�0i��A�+"���Q�;�ťd�;����|�&���Zk�����������o�w<>[�D�mFd���Q����-��cdhg0�ZP�i�ȊV��ۧ�*�C��*9�C���C��>����S�9B�?������:�'�Ì˿��n��?;?dI���3u�z�V1���m~�j���t�ғ�G����jkZ7U���~��~��~�H�^��z^����5���� ���*�"f~��,�.��3�5����;��~y�+M�q���2��!�F�2�����#L �����&��/&X���=!��ҋ�E�.}y��jzT~=K���I�yh�����P�p�hFExrj�6�8��]-��y��F�%��0��t'"��8B�X�lK=� �Ė��׻Y"��L�ƽ2�R�����(
�r��o1�<��$;��1��̕�.`����{��F7���ű�	��I�q�n��]�3,�v�}˶�4SJ7D��t~l�2�g�sXF� 2"<' ��4p=��s>�l�-+��D�_N�o-z�7��N�N�!�ͻ����q~�޽����0�<�g>��{��	��C�p����'��4���_ƅ��u�+�<���Q�⪎���F% ��oz�u�yiׄ�
�g)U��f0̱�q7�^�Qa��9�ڍ䭏�b.*��< #��n�f��]���}�<S)J �y�$!�x��Tr�#�u��]>�竹Auԥ�:9��D_��'���F�r����=�j���O{@��sx�PZ���龛�V��3��汴��N�"����»H�b��<їT����c��?U
���'����Xlҟ�0�զ��fY�@uDK���U�a�����+�� �uAA��Ћ��V*���ZBE����h�Mu�t��R΃d�Ղ���t�r�cPJ|�r#�:�wD�C&�-'+ o��
�]���$��+�"?&�Ѥ��@���ZF��h� L��,�i�٩�RͶRZ���������d)$�q<�i£+ �Uq�� ���?Ȣ �z�i���2��bcT����D"y؇w�f?�k���rGK*P���$hW"dĴ��8�Zњ�-|����L�� �D��u�e��@S�y �J=��ES��dh���ZI_ 6�Y��Z=��?pu��0;��:n^�f�ݛ���t�_uѶ7����gH`�?��M��N�G�����Ƈk�}`%�1R�[��%���,�-�ρvN.@1��/M���}���׍�m�6�,YKry%β�[�C�!�fa�P'l#������@>�cڲxEl�����𻲩�-��Ե�L-�.
��t�Vۦ��M�����<��QF�6�V&���7�O�Y�&�{�)2[�	ץ6�����Y�I�^�F)���粡��;
.H���a&n��]��R��hիܺ�4��U�؆�ye��|*�GB�m�-˜(�����O�2NV+�/Q�S&$�z9#��zL>�}�h�o������-]��=��ݚ���9d}QN������'�.����!?�D_��� j�����z'��~ϫ5���- `��_��$��導u��j�b�t��W�vHm/�A�afH�}�!�l����sﳁ�[��:������i9��"�� ��r��y���o��1I�ڼ��+��ctxd3���:���>~��jf�c�w:I}��N%V!�+�:gR]7�J�yR]_�d���rY:^������v'��)����)r	g�u���R2ZC���h�+#�?�P���E ��=a�յ��7쫁M�kD�����A��ş�*��[<M�R0H���zѻ��%p;-y_ό2j͋k#Q�}����b��
2���"[�԰�io� Z	e7z�Wn��}��u�Ocu�1�dq�b����,vFynD!􋦚��7�'�o4<�]�x��~'��� ;$�ȣ.��`��Kv�)�Ͳ�=�l�	tY��m�����|T>:�0|�f|:&�d���Kt&�j{- ��n��ɍ}	q��r5/k�o$��*��ҿ�C1$.�6D	�wY'͆�&���P-?�׹%���t?�q�����J_G<t �]��"䆏�x�8�P�<�����R���B�љV�:r	Lcn@*8X�t1�0���9�+h���AR�'9`<���Y��*����}	l/RLO�ֈ�^��D+���6Rjah��V����(�Ķ��'����z�ƛ�o���u��/.�a�`Sy��d>z7*�!�nA�-�.�����x��q��/IV!W3(}���_\����&�6��4ҭHD��h]�bS�m�w�C����k�x�l0s�B��q����ָ��
T_@��|��=�Ov�4sL �I��hW��P��G l>��`�]	cz\�P�|k׃���F����>�#o��M��.{n%�=���8bڿ������^��+�j=�����;R��I|B�.�^K��y��N_�̼�躽0sl2�2;��
!�����ZZv� f�����p$D�@�e��-ƯL��s�Ke��S(A��	8�n�9��E3g��{جc��EH�si�9*��h(�	w"y2��Qi
���aqu0G��%��*�B-YA[�P��#-�@�!H"�6�gx�旇>�g���<(��	cG@�.t�����ZY7@Y4�e�f����<q�ͩ�9�4$����}r0��t�k��>������_��ޛܯ��+�	���f[���}`���q�oib�h>K\c)�����-��o��r�c.�8��W�9��u����CN�(A���~��bᑀ�������S�T"GR3�r��tǛ��n<�L.������qr��C��J�o��ts	B����;*��f���+;�P��8���o����{�/���|p��΀��}';*0z3~x:7|��G�J�:�Е�.@�O8�o�{�9z�WF���T����ub�W΅�����Y�@����5
�<oAt�x��~���X�~3�%.��W� �x à ;����C�4%�c�� |�����A�Gmw2�p�PW �" �4�R(;��=#e����:���.�Ǉ3���
�2�镁m���2��F��j������>=�����:1����4��t�i2ꓛQ���|%X#�~H�J�C������d��lXh���~5�{I�3��շe�|��򼹎Iƶ��.��e����!������N�>%ĂDUذ�P�*^��^o'�XY�j6��y��Q����Yf��
�G���
��i��O��(�W�}�pP�R%���X�+�a�&����+�+�r�'��DK$8�9ýaQ=�HƢ�ͮ_��ׄ�@u� *���Ե����F��du5M�h��ɒ	Y!A�9JE-]�v��Va^xE5=>���K�	�t<�?c�y
��+.o^(΄&μD�X}l��1Ƙsyi�g���P�m�8��hz�9+�T��Z곁���ye���-b!���U�܂��<}�t��L(�ߪu?��vN5M�4��G5c����~��C�
?�~1�cIG�p �
�Ҏw��rH������Y�*#�
��&�S�V.L ��d^�x�)���3�g��d��:N?)�'�G�U}\��׼����奉��+C�Ψ������#�"�ĎZ�<s1<	gz�\�m��؀g���x��̯~=K�	APGL'}���1��H��ޭ�P���8 j\9��;�,=�/y�3Gc�� g!;rα�X��_�f������Kx�ܶ]����'�Ɛ���S��]8c��Ȫ�
����݅���>����\���/˦�H�c:d�Jd�:��'���87��۠"��8�5��
�{���1U��z���0����#[�ʊw_���Nqmf�t��9�?O!�o�y�TS�$V���oǱ�t+l�f�A�qm�ֹf^�Q�%W�� ���tbsBe�׺�jd��^���H������>�i���/��ڞ�ȁh��*� ˟�$����M~��W����r炊�_iE���:;� �\��/����M9&�̮п&�^RDI�|HM�s�uq�#�c�#PG�p�"��J}"��j�lN�k���{z�e�����BDB��EJ�e��� �7��*�a4�J˒^����~��/VVˆ�Fk�QhGm#-\N�ӿ׍�������=�u�C-J3���'P��S�u���䱨-#�^�`�}�Rߵ-��P =�}���������V��k���N�*;�A���5�]�7ފA
A�٠��X�sa���0�o ��|�	,zCF/b����U����$��͔ 亵��&I&���a^���{DI�������J�i��t$�P��>�����?w���V���T��밈au�v���MW���rm�EФ�ܟ��<vςS�Q)�7�ɚc�*�j�]��>��L,L�ڑ�Y�+�Brp�_1-ˀY��&�A����2��w��%� �1����VvN��߅���>GH��K��R-%(������u�r�x⏎!���+�	��K젂�Ң	W�Mr�e���EK��qW�"��M[�$'5Jj��6z
��P�^fv ��iJ�}�&�@��t��	 ����JCp���٠,��7q�E7���f]�{��-:�P�v���,��U�Ltc�������g��S1�=��Qb���dҡ�8��2��m��k��T��g�p��G�_�ς�k�ИՃ9M��nL� ��dݘ����B��/�|qDu r��;���c�r��=xw��e�a��܆i�8�np�S�u��0�]4?���ɽ��k,Oa:p���3��
 ��E_0�ǃ?�n�����b�gN�l�W�8M;��&��ɣ&�1�l�!�~&{wT�l�r2[�g~ح��[g���B?�����w�F��byѤI.:G�$H��9��_h������IC��e�i�<b����I��{��U8`�6���b?#'���8�f(�����^G�^O�Jƀ�����{���D���d��(�'�j��7�X���$���vo�Y��p�]!*s�H����T�A������p��(�}[ֿ��x����=pGH�Q?��2��n�A� z�W�����iG�G�Tg2��G�
��-�5Ř@��L�e�s¥���H�W�37Tg�{RY��N��������5~�@����?�XW�k1؂E����'��� J�:a��4bh�?��Z�i'��m�"�i���έ�T�H�%m��� \;J�X՜Ke1���M��������Κ~������į�U��C�ސ�+���Z
����g�7?M)D�)��;J�g~�H;�p��c�}v*{r�|�z8b�m�G^����|yRni'\0��^�f�_�vS��)��5�f����|`�e��b�����EKb�e4�L���v�|$b#�=��M�C�Ѵ�K��,�����x�#X 7��q�f�hMY2�Bx�}jb-�,9�:Ej�Z��%Œҕ�8ɕ>�Ӕ5��_00�'��pbW���G����o'�\����z�j��C'_ ��k��z�?V��@�'�]tW����M�P�Tc[v)w�t��@���-�y@k|���'kֽ�	ic����>��*�Pc�Ü�^.o7�m:E�`Eym�o'����]����|;�-��]S��',�|ĥ�@n�;$��w�������C"��k����BU��	�ؘOSX�.&�g�儅�Y�(�h�>���2�Bf;����54X�
�0,o���n�C2�3gn���_�y%y�`��E�Sl��"1���ѥ�RQ��;��<�c���h�8R���+\>��c�7�j%��nG����9��`��4�XlxVHYEB    8e10    18e0N�����D��Y�V�x$:��,��v��������4�3jY���-�5M��[,�D:��RLUָD֡2��ǪzZ󔧰�܆���F�F���9z��_�
��Wa�!>(ћk���gH�&���{��~s�X}��+�̰��_�e�b��2�@���[�ZY�܏�j�,$��7Dm�Qk�ϡ`�)w��S%���3le,��*&�( ����4������k~�p{[����,�Bw���n�$��:�m���mӫ�OVN�K����;��r�^�&4X��|��d-��淋I��H��1��ڔj��.p��8P��1dU����6�/� S.���L��A�Z�����E���B�[�{�x�j Ԗ�V�� �V�]�8Lc���|�ǉj$][!�F�e���2�m)#��@ "�|ӟ��3�;�D����6�ʃ��Ĺ'E����ɶ���Σƹ�zQ�t�Ai>}�>ێ������.�R�÷�2q�Dg����ߝ&y�O�)�����X�A��Fav�%^O�M@�;���hheȦ�8��R=k���{l��  ƹ��w�r���[������p�g��U$��3�D�xT�Z��C�r�)��[E��H��pۛ�:���y1��C�wr⏻V�9���%V@pԖ%�HAk�P�\+vaL $>}uUE+稜��l�����# |t~&em/����!2��T{m�<��7{�"�<��v�/�L�U�i��3�'����ڮ|{bJ3�%�����;O�	f��;��Z\+�܏�x�5<0�l�L�PXѡ�"Q�A��&ș�c-�����-�	�6���8�tA�F�����[-�F�;�$���n�Fjen�g���ޥ�Iu-�ezp�AKBFSTh��΍�FH��q,`C�L�uD���eX(6�'�BN�,��e�|~���j�6Y,��n�!���׀ݤ%�V�"N����QV����"��0t��%e�}j-�o�X1���y����(m�ÕI�a����et�}<�A,���D�zN�A��4�-������p�ں.���q����g{j��;���v�k����tx�ֺRPt'-�OEԗe��~��aC�gpW�V#b�'�ǟgD���Ӌ�fp�g�P�6l�mXvw��L��7��O�)���B��� C�=&,\AK�#�O7e��趜��Y��`�3&q���������<,{�Ҿ��n~��_��]xHH<l��ϣ��#x���Q4�>��i�^�:w����$�K�+�$�u�;l���i�:�P�/�
/le���~^)E�t���e�11A RT"��,�t�G���~�a�$��!�F=ж��$I� �j�s"�̞���^���P���G=P��X�H^EV	�ж{�gv��G�G���n}�Bn#��g��z��[[�����I��t���kd����GU�cG��
x�r N*+��r�s{�za�$���E��OQ@y�$����S�q����jZ<Q�aӪ���;�/�M�{�P��`H�ff��9�<c^Nt�ta��J��^��ki��T5��q �>"�FU����$���<����������P��)�f�iּ�����0�9��vdZ���S�S�
X~��m@��S�oo�s�GD�`��F��9�U ��Tx�y/c� �ՈDq�̀��$�Bq Ě	�)���KK6��hb��L'����>+�w�=�w��HX5:y�����!YB[�����/u@�]��y��:?Q��1$�B��C�2����lE�}s�|瘗������w���,��|s`G�`VU�~+Ѡb���%��k�̯��
3��G�(�R@v�g�ѩ�V(k��n磙��������%�ZY�!���N�D!V�0���2p ��T��KX�`�u�'}W���@`��lE�^թٔW�a{��Qy�a(G��7�lQ��:?hˠ$ԃ�C��O&RAZe��6���%�`e�X�!,��rҏS��:���P��w�{*�9�lҾ�n�LPF��:�Y��Á	&L��07��U"��y�ύ�ƻ<�?�
���U^X�zr�D����9������{���@ YA�xĦ�%s�F�Gas����m��v��s��:���
^*�nKf��̞�o�{?*%v�Q� �P�jvUs2�^�����f��s���ɺyny����g�v�\��nQZ�͡m�R~:9�I�=)d��\�,���Z
UG�6��I��f_�jѸ��i���&�,4Cir)+����ǉ9�}�`B�A��l���C6v����<�V�NE:�߇i��9��]�CksD����Ҡc��*���}h26^�V�bT���$fb���M�f���J�o5��
�,1>q�8<���<o�ZJ�՝�X$He���k�z�f�!J���g/�����B�Λwq� 0M�|Ry�=�$��=�<�Ͽ�}=cY����*�� �ɿ��Vך��~��/���&���^�ɑa&��Fw�.�_ҁTL�.?���]���lh�"��8n����_T�Y/� �'�[��)*���;��i.�c���F�]%M�*��@U�-�
�wsމ�n$9'紭�-fkA$,��~�NO\cii�v�E͙?���w�qrmc����HL-�̏!B`�5��>���%(p/ �Xc5�,�o=uX��n�d�W����������CC��`�nR��H98�#�5C�-H�6v�% �:9yQ(*�߇��,�*]B'�ya&��Q��DZ,<�ٯ����?΄�:������#t�-�=���0�\���/��Y��*[��J�ߧ�L�^{#�l�}��>����˸	�8���f�+�o�Wā^�G�|T��ϯS�}
�Z�u���j>�󊘅��YJi��n.B���2%F���7��7�m�O�Y��
u\c��Ep��i��c=Z��@�������h�4`n|��:-�έe'1�Yw�L �bp��b��h��<�W�z)�OL���3�2��qӯd��T(n��O��k2��x��m�2�ƕY�gw8�ϱ���1�8"������N��ڤ�@�f��x�Ë�k)*�����}��~�'l)CC?���x=[V�[�[�_ ��U�9��rG����
@&�����ksa��b�"��� ��d��8�R}�R���
�k?��!#s��,��C�р#�/Ie׃����{��n��\���k���a������5��4.h�b��y����.���O�(L���������mn���m0�J���	+ţV'�yXE�tŢw��QX!;�2j��x���1�}��^���Nܮ�9k�8��r��#����_�Ą�X����_j�"zՀ����i�J�>	Og���#:�$OR��u�\�cwqE����퍬�j�d�&mp���U|�PngPn��aSɟ����`�iycn��O�I3*K�w\}�i�c�AviAXBM<H��őa�A���u>A�G�ZH.N�J4�����Mz�ZXP��'dF�?+Y�ñke�
�b��A�U��WܩD�Tދ~�Fk	���I ۼ/ɶ���
�A�����9�2�XD��� �����/�p��0:�.=8�9���40��vdbܵX:Z��:K[�iԃA���p�� o��|c���I���&���2^s��9Գ�:`�����-�ͷ��gZ2�C*�I���Ӏn��3N�_������cu�nF�1������^
����5;�$	��+�]x��&S��z;�4D������8�2K}v�g�ސXX�������Q�$��a�n1q��zhu��RY��I]}4u:�wibI����.ٯ����|���a��R=#�����vRqJq��E�58ߡs���l��i�f��󌐱������I$��E�I?�!b����v�/]�)`��n�64߮/�3)ީ���=I�߯�72�|1�Ki���n
�CJ�����t'�?5=6N� ?���� �];Nj_S�T�k�(8�bR�)=��V���@k���qq���y�!<���d�8RҴK��C��Nkk�X�ޞؒkL'�ӊ�t;:� 0Y��ٜ�f۬"vͺjqidUu��T�'��P��r!LltG�4hŒ���b�| ׾De	Md=dތ��N%U�L�<j�4�\�E�F
�p��?������Ł���3),2���i߳IA�?�m.���s���JJ�Җ�[�m5|���64�u�6|�f��FҚ��<��SW�8e�o�`���kq�[��5����a��һ�W%�i �'A;]���P)���IQ�e��uع-#pL����׀�<�g�$�ID�0���^Ѳ�'�c:q&nL�`:����r3����~m��\�:O\�~���D�x��1	GjަC">�Ǵ��2-� 9i�_���������j�Z���^k���ɺ���cMb�Zuyx݅��S�6��Y�\�VB[Px�)�:�tv~����O���*�ﴸr�}8*\�,��>�i�
�%�xe^��s�r0���y^ȪK�br!��ᘍ���q�\�Q��������4�@�@aP�IY7�л��z(\��W�����Db͉:	��Y^��q����;,�ɕD@�tӁ�0���W�?ۮ���8�t��\��IY�`��-@�ϯ���!Cj}�$V[@+����iYM�z��_F=G~�*��o�B�ŝ��fƔ$E7�in�,��#$}j�c� Kb<�p8�OnY�>��kj����l�z�)�6�����}�)e����9��<Ǽ/m��i�׹�V'���s�,[>.u���j�dE.t|Ή��E@v�������1ތ��0G�3���|��������h��<_���̑���Ra�P�9m@��\X�SGu<�æj��JD:���M%qJ��w$�wjD:��v�8C曃��4��R:�!'����3=�L��2�c�>�8���[؏��d�S����ނ]���m�A�M5�r[Ɓ�$�B7�YD*.�x�3�1�U!M(�?���08�(�=q'�|y*9��Ae�Z��<�k�3�Q��X�Go�%j�$����,�"sbb�$�Z~�c'���zv�~tby)k���(so��O�U���xR��D�k��2�D����Bv��}?�V�}
�>`�(����! ��#�I���}��ޢ�t�U���.�w� 6 ���o�'�քpx�B��g�#�dYܸ� ��.`3�� �`L�=�-�u�$z�,�N��g�C]�nsw�H#��(�W:X́ȋ=f��wo�6[��!;!��	�A�-<�JL0�~�ѣo۴@Z�V��}��eM�I*�	)i�yvN���6-P�+�-��[$>�ަ�K��-�r�kV��;��*,Փf�yn��}}��qIA�9m�����:��h3����đ~�ɢh��+�/�r�wfFZE���|\b��J=8m��4M6���_��|��pr0gd����`	�#�V�5w�a��orM,+7 �_��5H�
v�ծé݂��j{����^q�!�(^
�����6`�Ŧ�d�lT�=����GEMh3JJ��$�f�Z���؅����W_5����;:��x��/�R��Yj��{E�l�Hh�m/o6���FF��փ�����v�dkA��蔒�������c�_#,��I�X�:��Upk"?�����~$�J���{L`Ó�!m��Q����?����_�f)���S��n�����3P�Q�o�!�Q����0~-Rktʠ%)�
m%����i�G?!�7��FQ����˴�i0��OƷ���T'���L,��p�J�B�(�q֢6����c���r�
TKx�:��i�c�JF�M�?d��{9�t0�Ba�&_�Ϥ���?�t��^4�b�*Qw�x)N�۞y��0�o�&O�kG����p~�����;'�����`/Qdׂ�����\Rݓ=}�`��k8�TD��QǄ.'ņ��lq剺�&YJ��K�3�50���eN�#�k4E�Чr� Lc,+�ۗ�d�ϊ��%jb״��&�f^)�I���L����4�f]c�/�����=�hs�W���m��y��Xp=(5��{�B=�+9�O��a��K�p�Z����H�R�v�^[)�dsQ#_��F!�\�Ĳ�(�$��v��۵��R`ys������^8h���)a�G&���p|���g���jI礋I�K�