XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���̿C6
4�o P�{r��_��{�P&p�`�D;=����S�?�5D����w�M�n�QC�'��Mc���1 7{�d ++Fl��9w� ݨwoC��@�X���3'�U)�������Z���D�N	�r!J��/T�ipY�нJ)PN�*�9y�_&1$˕)���+��(@��X�����;ӳ ��AgS��>x�����v	�5ج�=�a��5�WiDlZ{J&f&�W;u �4�	�lx}_@H�|���4�2�*e�7nK�k�����a�f�$�H/)�4��]�ZF��sI���q��8���z�&7�G�_��������5��!_�r��X����H�H��sXw��N�u:�U~.�x8A�)\YL�d�'2w����?��1��j,��=�/��Ev����*ƫe^z��]Cu��.f�AF�HFES{bq�'Iԓ�Tj�a��U2?�t߶�������8�'��	�E���aj�aG��y+��8c��tgw�dL����SKRܽ���NQ��<Sge�IQ�[V��$Ou��P� }C��F �_T�we��@e	��p	:<��)'�q-�h���[Nn���ᨨY� �g�� ��_���B��ࡸv�\]bt٭�p��(��MsR�-f��͟K}��Y�-�$��K�Tē����z��� �f2�.lr�c��P(&Q�ܻb����G����Ug�R�U�!�"c��]^��Kn)���DZK-ǁ2�>
���.e~�!��1�XlxVHYEB    fa00    3000��r� �A�O�D���T?rL�5�+��^yl���]�Ϧ��J5f'���#�8����y��7�kԃP�)���-݆{ϻy�`;�y��h��`�ǚ�uƾ�b�̱x*[������!�,��?�g��Au�I%i!�*��	�cNB��@-5@������+��\��3.&��c��(�4�f4�B����W�Q�g?Վh�׀��G�佪E�Ҷ��Q �"&����ؙ��|'�o�?��s're`��8��Vx�P1��I���	�&����g6�o �o�#�Wfa��mTA��L�,]����������矄�1e�a�q�`�%F8�WF�%	�3�{/���"tӤ_�hd`�:D�ZrӶ�>���l�Tl�u�u��kϞnt�Ә�T�&z���EC�A��]��yLjt{��_�@��,�8�L�k|p��?��6�)���˴�;��e"��m��c�u[	��A�J�{ᅷ��Q���Ewz`Zw��~������(A�8DX�	�[�>���l�k��g1�/�DA�cG�-��7xF�y�x���'�=U�TӮo&���k���j9T���ܪ���53����<_�X���T?�"ŎA4O��`��j *����uԠ&E"��D�mx]F��g�峿o��?��!�O@�!�Xp��q�������E(%�	��H��Dn��*PЕއ}���=�~��|��!�Rg!A�~P~��<�&��� %6	2L���!	N�'|�{�����TMXo5tR�%��P�뢤�2cP�	9`-IlE��iܕ��J�������G�V�@l>ܸ�I?{�$�P`��+Xf�y'�Z��{��t#|����ϻ��ؠ�lPد���Eԍ�m���#��Z�X�[0l�3����C@��hXx�f�d}6ۉ%7�\8'�������a�xQ%�}-�IS�4%���+�"4�'ä���+�ҋ��:���>v�Xz�����P�콺�P�����"&����6	��� � ]���#.�A?�����D�Z�n���
���K�Aq�:H�y���n'���)fb�e^5��z�B���j�z�:�cBG����)mG�W۵K�y:�U�0\�":Y-eN��e+o�~�!n����ikϷ<m��)�S$Ꚓt**JG��/..�}�bK\ܽ���[q�#jZ�?�#��Tn*�������O�X ���c���8#۱=�����_�rP<���_�����ʪѥ��ʷ'4R�)x�*A6��7�"��Xփ���4���D zw�8V-��	��\F=���L����7�8���a�ԳK#�s�Ɔl�?�83�̾jo
���k��#aZ�)��gz��@����:�##e� =@8)C�[-�l�X��z_:�yR�̓y�R~F��+q��{%@�m9QͲ͌��t�̫�<�$�|S�_L	b)fU�a�n,`�~��afz�R���*�9�+�iF��FъP��4؈��r�L�?�e�0+;<���z��h�'�KA3�ȶIw�{��ʰH���1�;$W�5
h�u�H��S`�;A����o�[Q���Zq��/k�Gp+��P���@X�D|d�{*�����C������ځ�~VH�}�HP�?�Hֻ�An`��v/
��J�ޒķ|X敯'��A�)8_5KL�5� ��N^�����ę�N]x�LR���M��U ��f�{��65I�g��'���]#p�X�cz~���:�Ǽ���+��O���rl=o��o���>�ԁ�Ξ�=dc}z��	g+��jkW���	�E�β�m��f?C�!���te^������k2�Ⱥ������Ot����wt��yC�#䄵�`y�����9�+��By^F(�)��á$s�a#u�1҇�g|�����P��$��*�)ti>_^6�УTvG�������kjw���$A��o�F�ڭB�?�{Gl��>b��j��B��W},�h� S.JO�ؐ�D ��4̏W�A���GZښ�M5�!��Շ8��MS}������e}�p�ݙAG�i���v3��!�u�/X��x�����C*"�߈��=>�J �]r*���2�
�kH�栐Dq���������0߻��֮DF�h)��2��>����TY���VP�� ��i����t�Nίe	����W�BJ0���P�d����e�ε�\�� ސ�� ��kp9�T��j}�f��S!����Ie�H�����3EH��p+�G�ɛG)A7��qc�w�n:���_�KW |#��.��ѷ�:.({.��d�y���v����~�R͵�ē�~��E���5����-k2�<*3~���GMY�'L32��VR�����+c��B�{��3��4�|�PЮji����z<\tu�����̚��Q� gl,���[g��a���?`> �4�Z1ۏi��pؐ���5�Q���W��'���0(�b$kO����T
�-Q9��c���y"��D �@$��R�=S�?�=�K�ݝ*e�Qֳ詬����m��]p8���:n�_O%z��AQO6��$���2����L��sȡK!꣸`L�Ци�V�X���Jq�����h ����Lo4&3�̂�� �q8cq���rUh�%����I�k�S9Kr�[��O�Z��Y����5y�5�ms�5S|ݠz9�2��ΘB(ƽ���S����\�t�9+	I�e�j��n�ߑ8��}�|z�ꍑ���^�^�G��+��M ��\�O+�T�E�e�$[� sԛ"k�^����P�����.-��s��ː��ŋ�����%�}r=w��'#.�)��Q�1`��x��{3$��������-/�WA�qTE9�������NS���I��f'�%l=)p�^tST���z�V?����Y�������YFKzTt���X�g���]��l}���"��ޔc���L3O7�g|���]#�X�����C .�j1m�I�r������R�Q>5yv���9Fl	zٰ�'kC��Ǔp�Ju��s��ix���%��V@z�)G'��!�jA?�*��X���,��
�E$��'�+Iēq�3���ft'�vc���nf�4���8I���$i���^aӈ��	W�V�6/�y�z��?��E.��n}* H��
P��CB�� p�8�I2i��-�0�����O+m�_Z@�<��Ԟ�!h�Ǘ}�B`Čh̝������>_�n��;w�f#Baĉ�ħa����]h�&��A�gA�FD�@e����#��H�*�.�Bh�X�����k�p.Q�j�0Q��]ܞk)|ڈt	�Ƞ7�x�T�z�-��߼�V. i�`"�IC�r��hu/{d���l�t�!������f��L_���?�����"ٸ���OyCO|��.\�&�~����A��x��jp�
��v!�u����!�H��!Η�\@}�?דsT����)r����DN�-ʴ��C=�`F���|a)8�MP�x%�]hg�}!�ȸ����b4�>��>s�=Y�:���!!�ܔW#볍�E������[m��@�R�r��P�����ʞ��H�hR�Y-� /��ė�t=M��v��-�YCi������6�I�����mH��N91��#餃j�'�Hq�d�7M��۵�i8V��y��h�7�{(�(�&t!��}�b+�o�W�U�0�"!EM9TwV�H��>�XZS�ysEgcp$�	H
قs>Ne7^��2<C�t,�;�Np�2�LJ��q���Է\D������n"���]�'P����k�g���=��,<�2��T鲕\�D�7�J����̦q9*�tH�T��ְB�	T�z?�J����.�<�c���4��ڂ����^0n������P�Ni��Y��4m�RӺ��jK��r��v�.� I��~��5�ʗh5�j��Kr<L�Y�u�^��MF8�2\���ͤ���1^�r�������E��s�L��W�~�=u�?i��	�ӥA�8�"^>��4F:R�mD�S�I��-�X�`�Ú���1IM�.��)l���mǼ᝽��s3���$��ކ2��С��;�E�'����=bf��&�d���aڳL0aNt΃�pG���,f���)�����OE���ܨ�C��~�!^W=�O����r�|2@P����'�}�]�����:.�z�O���P^]u���!���%�7&�T�������t.`��T�1y�j0����nL'�Ɣ<=�*����ck�ij���ȧ�A|YAq�U�OLx�^�8��L�:!bg|�e�<��IqV��7�M�lt����倯�bko�7�z-���n���Y����7|L1����+C��8�"���;L�s�N�o��U��u���+��Ty@;�3 z6��Cv��^��}H�5	a��u�J���=�<�x�;҂�!�	o� ���Q���$�7(�'Ɇ����^��z��~#b0����;#���-��M�T��fM z�t���^N<V�Q�����2�����C?���ْ��b����_4s JF�ɼC��kN{,�ng@���q��*[�<!���f�v��rӖPnMd�#En��T��Ś�y�ןN2�x��HgV���0"ѲΔ�/v�
jJ�AE_ ��(�����~L�b���g����ໍ��g�S]���J�3*�n�xrhaZT	FCG�{��0~L�=���p=7n�u;�9C�
�)7��!�*����~Ol��q@�Q��W|_��������3-����_As���_�n<~��K	�io��e��C���j �} ����߄�?�Q���8�Ld[&+`��g������7@_�Cݎ�{�� l>�Ab+�,�8�rD���Q�G������Zs��jy�S}j<��7�+1��Fy�y{�w9���Cn�gQ� �cEn��l��a��m��9a%"rY�
u�1P��΄$pk���y�λu�%���L�*���%.�D9+���3
>��Xⷉ���[a�)�oW�\�r��Yr����R���?!/��Ch�^�b~��p��Of%�j��*������~�"pW���W�}��i"��;2W��Usp�i1ܬYk8��1�a��FC�o�B	�$��Wwr��DsR�����Ǻ�"��1��q����
����
��J����'�:Hg�x�m-����m��e�Y vm<�S��m�/f�k�5s�.t��0��]t0i���&9G4!{<�Pqs8��� |L�b
U��^���=.Y۪%$5�V�R�H�*,�>F���R}ǟ&�C�l۝�-��/���^A�#�p��曉qC���߃(�k��dۆtk�"a�A�&Jp?r�S^b�/r.X�bd%�睊���S��Y��A5G^:��@G�t��>��z�
�^��p({���ț�r�m}��u=�!pzP��յ��HY�8	(�%�qv�'~��l��F��tG�P�q�i�F��E�<r�L����8>�ةN��R㚉c�߼��{r�,��f�P�GO�&�uT��V�&gx��Gfū��:7������?$��ԓ�X�����-�F�XQ��o�-��
����.���ԓ�t]�� D0�����z�]���$�'�6���u�<��~��[����@k��ߥ����y5.��L����h��k -�a^T�09"�ЌG|�Ő_	�'�n�u�Ѿ*��ă�!aiGz���%-�^�/b��c����UH���^��>���z�;\^��k�kb����U�}NDW�K��~|���{�p�����2�ȱXoܕ+�	���8Nd�>��^�ԇ��?A�AD���ٺ��=��d`V��A�[?'��g�y���Q�L{��."�N�b_��`nV����Ik_8�>Y�eY�m�׫p�q����Ǖ25̮���k&�m����#����l��v���1w='�*���X���Д�����dbZ��m�4f\�ge(J�^LS6��V�t��z_��[׺In���Mɽ�<�RM�/�?_=��pNEvوx�zW���C���En>��_ŎJD���ʷ��=+oҡ|�Ϛk_k����=R���a�ـo-K3���џ��1���9?���z�J���yC�$�c����E�;�T�	�6n�\�M�̢���?Ƭ1I��C--W�7S�^����N����0{��M'�e?y� ���0�-'���kcMu�Ͱ�F����(Te@0�]�a^}�glvX�`�t�SB�8n9��\ Ze�3��w=@Ǭ�lø&?�ftc֥��S,CW�ȫ�[��@g�9�!U��b��۱��t�֢�{�K�dr�AiGO�lx�1{�q���7d��s�s�p%����a�򹌟?�9a��kۭq�,�3��>zye�1�[WҤr)/$1A��~����ؾ��6�W҂��rSI�SX�DF'���`ş����U�V���=��Z�aj��I
��P2>"n�qT*:L�
�Cy�{ai�ԯ�����y�>n	GzI�kI7V��xD���*���3g��ޭ�Rg2��v*cv�=qx!��@@���#P5�ίT����M��������@�%(���>`,��к����u�kz� �E�M/?߬�#�nӛ~r�p��7�XGf֝l����=�<s�}����2��ܮA����Y�Sg����Ҿ��[�l�|o�ƛS�1�[��:���#��&�nR$)�us��xe+Q���C<����l $zh����&:R3kG��Mm�ؙL�|����)�H�
�U,d�������޸�v@z�:��8&��o ?XA.���P�\�0�/7�,00���=�#��i��2�]��O��ۛ�Noriչ�i
A��"��F/�kƿ�3�����BLjւ:�������T��~2��ʩk����Q(�p}��}�T�w~�D�{U��*�@�6e� ��V�~�ņ*_	�+Qf'j-Q{f"�eZClq�~��Qm�49x�,a���nN譢�X����?�t�ef�W@�0��d��p�Q�����W����н�BW�Or��h�*�V������Y�4r�}�Z+�qXK �����E�&�h,	�?t�2:	B,�mb�5��KJ�`O?X�y����xҡX�۫��(N��э^��w9����n/�M6[-�;1��m(�	�7^�s��t�J;:����"���͸����ۚW��S����i�ڴ[B��M_5��)�!!~�RҤ�����Yy i���ݝi�
�#�V'�V9������n
2���+�����dg0�~潚��Vև����%D�mh$�rG�FB��ܛ���\4�����dG;�3]ǯ/��2�<n��x)R������?D�=�o��6���!���X:��t	&l�`g}�b>5�Gպ�օ:r��-��I�J�����r��6	!�8j�;��=&��3�u]��}��evp���ߚ� -
��ڏcs���km0J�@�����l=����2��4�Pٵ��f��A�����\85�ޥ�F-�֒���G8�µ9�$�ͿZ�7�F��a��n_����"B�#ב���7��e�Ά{��^݅�//�C-,M�{���Թ��B�"�QϵC䶫O�����:��vx(�U�/�".�����k�/n�ZCߢ#�
�t�n�����sO�m3��4�V��\���G��B ݆'�l.�h�P0R�L�!�ҶAE.��yC����*(ei3�1�^,�ps�ު�#�>�g�PX)�U�g�R�S�r�S�����q��7Ӳ�T"Eo~❷��=�9U���A���E��DAJ#^Cz�-�=��<Ӆ8�R�^N3@ȮQj4����K�2XA^jϏ�|�eܝ�x���i�X��&w;~� =��73��9����Zq��z�{�S̊�R� ���y�~��+y�C.3>��
y
>o�@Y��_����e#k��N]�w-�{���#l�a/9�+�Ϳ�>�\ƥ��ͤ)�,�c����d����)A�^����Jڿ��ǭ[!"��R��ˋ�ւ+�)�����.��Kڎ��o!S����+Ӽ����;j������E3w�%6�ݏ�Z%�1��r��J ���J�$&"Ň�������c\��{`׶t)j�#
�m�6/�;� ���D���s�lin���b�S��!N)	fIsk?aZ�WɽŽ����8�b��/N��C
�х�ֽ/`�������0s|���ڊ}���>�7�/���_�y�/[C3h�l4Ap�����^2Jr�p;5��v�{����J�!	N������JE�Yko~��@�{>�M5�ϻ�Ȋ=2`��ڙ�,m���?�(�n���j�o*ީH�4��	h�;ء���.3�~Y��]�Mu���|�}��ރ��%?�� �&��+��ў��{	�|Fn��־��O|������{7#9��K��B�a�j>�z������
v3���E�������f��R#��(����#����E��1���~v��	j%�}�|�=�ނ�h�*�l��z��rbu�z������}��νE��2Q�seT����ɯɾ�rWW%����	��g��������I;��<��ܚ޵c 
����5d��~;�����Q�;nM�s~����0�c:�^�j��B��{!��]:��j�����WK�9�K��dF��ݥ_��iH�������7��:Ib(��[.S�L[t<��%�M�j�W��Q��I��i�cl�-��(V��c�(����]_�Q]""�qo߸�x
X��ĈS1���g�.��6��|�ȴ���A�̑���9������k%(f;h`+��!頏�����Y��V�U�&{�=�����ZEC��EZ�Qқ?�c\�z���п=�'/�����+g�:qb/2"��<QoM�/���Oӡ0�P��D:�yj�M7kV����)C����FS�ꑰ{X8��ә,X�&iPR.��$'�fk�[�x-�^��٨���.�����l�bF^�����X3�']9`gL��v�jy����T�7r�O;vI\�Q���[¾-�*y^i��e��}$��v�}>�}���I>�#|�+	.qo2�
{�B�*�V"cl�-�6�D����D�B �g�ͫ�$<�<���g�>E̦9�e�e��oqk�:�����rK(��(���`u�sy������-U�C5��'A���9�S�Ě�,��Y0����i�@͎(!y+:K(�����{
?���{�_�p�T����<M� ��+i�7~�~>}�nOos(P�;��ۖ>�w:�+����z���!�Vo�	c>i�V��;�ݧ�8���`Nq`�k��E� >��e�3�E`�>-�_̢2O�yu�To�l=$8�%ϊ�'afޑ�*ԁ���4�z��QR�@ xJ�*�C(��KƽW�
Ϲbc�iD��&��Z H7tUpShD�`�/�����<�w/D�h>��!����B�:�>�6��9��
�p��T0�}F<��B+Y����hy0��I��7XL9��&�z�q��9؅#��f�h��21�C�6���#	���S�2�@ޓ�_z~�F��b�<�2]�	�x_�؃�@�~���Z+ ��cY4uwF�$h��ءT)u�������-s>B�e*�2��ޖ���q����l�Gc* "�[��Gr��9D�2Gc@R����s��3�	�s¶(��Ǉ��o-r������áȎ�4��V~�J?�;�c�x�oI��\��O;���p��\�����WG�s����~fȰyK��c���f2��6�]��d��(�ߎ�:�޻GO�̈+��)���Ԝ<f�2 JW��Xw���q�&3��u�E��}kB3�C)eSc�mi�[��A6. ���!�[5d�ɝ@)*cX�����������&����L����G\���U����ԛ�(]�."Cbv�s�L��7C������P�b>I0K>��*�� u����Nܾ�b"
��zi�������#֒����XA=H��IoN�6iiP�s35k �A�T��cH��;"<�)��n�Aˑv{�l���X��~�&��/�����[tT�|\�{n%����}6�-=G���N`���8�mNK���J���F�A�s��8����n��ҳ�>D�"�0�SxY�F����ܔ�E���9�|���)<�kK���{�����,p%�#�+��)U�M^�����YL�O�nQKe�޷�N�WM�)/O�	��)�ڼ�e�G��&�-�;�NT+*ѨLjcl%yt�'`Y��$?���}���L5���Q���#���5�w����dj��S����K���>4�6@"�) x���FJ ��y(�ᓠ�;�^�R�?W	���lSZ�4�r�-�w���C=�uQ#�~n��&�A�m\���R~���$�Gנ� o�.�YQ��l̋bG������b�	�� ^o4�tW>�D��?� 6B�S�%���'~�b�u�M}��^�gEP�}�K}2���\���Gg��T*�⟺�1�9��C�p4Qz��<L 'Aچ3�����@���{B�����}!�,�9x>�(j��޵��b|����	�_u�S����Z�t�~P��QѺ��3.�� 8��d	��x��MU^���֚�XB������<�]�ȫxJ";��Q������R�3�u�eԬ�Y��Y����������SF�Cn��pW<r���`&���R�e�����~<0�+�GL,�@��̨�3�Iޛw� ��!�A��{�!8��B��x.�NNPghE�UD`u��1HjYTQ�<ׯ����,xdri�k�9pK�g�|=��&��sGݩ���hg�_��Q�8�����T;���Ekgf��TF�D_�U��f�2�r��� �U��»�8�7*Wj_��%��^��Yg���G鲼Mx~���c�C_#.��Z���Y��xי6[o����ݯ��au+�U����$��`8ǂ���Sj��b��_����삩�ᛇ;U�6��ɑ��Z���F-����Vu���W���	�	�2^՗���L�C���[0K6̪�PŞ�9��W<� ��(������&j@�0��#y����n��0�1����F_D�0y��(�`�>m�TC�v;8J0M����OEJM�Mz'y��8R����M�+��U!N��t������X!�݉��4$�YGط�I~�ЕbY_��f=(�����qt��s�YskG�0��x�����7&��+IY�$��=1�����j�~�	7מEB��p�BK�M�p���W��������8���u��@�q��{�ܠ~��u~����o�B��о��?��6�U���d/�D���&b0�p��B�3c��?t���g�A̹EU�UΑ�Ԫxc�>� h��b���{#�Ag@r͠��9��g�M�;�ddr���3���q�jZ����~^��*:8�|y��J��wߊ�����G���r��o��5����o_�d5��X����sW|���R�yK*�,+����#&v>�F Ͱ�B��K�k�u��0��.<�=��S\��}
)��;0����`1_�]�=2��wBh��B�Ք�$�g+Lxnt9?D
v�J���)�o	F�>@��ROD)��-t�Kn���p��}������!|p�����������TA�F��ۆ����Y����ݓΏ�g��0j�����\�eR�;
�dx�0X�|Q��tC��"b��,`6Q�I ��St~��R�v�
�T����gC�/g8���#���̿���X�[1Q�c/=VQ�l	
$�]�( ���\	�|��b%\w-�;��{6W��<�e�i�s�rg[	�� ߍ#�Vl�C��B��:.h�W��F�h���m��̫�v[4	1����7��Dg�����&�ܹ�`|#�_w��f��Gҷ���+nV'��a�:m��y��"V���S��!ցK�]�Fݽ��6�#�؍	i)1�����#�f��XlxVHYEB    5ecd    1310Q4�����eK�N�P�3���
)��*���s~Q%��O�T�z�`S0M�Z9{a9�ωKʚ,'��Y4�E��i$�w�DrE�)l�}�.�7��������	������;��T�C{�+�k{ќ�;6D}��e1��n8V�������� F�R�� DƤ�`��\�i�P����Ɔ�&���8�-��$	�g�R��d�v#B�:���ta[A��;����F���bǰ{	�3ϔ9��=��=���8�n\�Ȑ�?�_+A(tTV�NT��IE�v����N�-�"Z� ��%�xκt6��� Q;K��������ec���BZ5����?�� �eM���z��z��=�����P�_<lM)Z��|�(���u�,�M�1L�q%�@1"��#���:���N��A�C�>�8#$���%�;����:m����k�z��t�AI���#<��:Ba�o������h�[�v�Dxm���j���Ʃ����6,6�y�P${-��7�{�#|SQ�#����wn���Q^��!��L�i܉,$�򕫴�]iAwLP�_���6���D,��JZ�&�U$~X#Q��3{@�h';�5ʧ�g�A 䫕�nT����Gu?Ď���{*|�����%ޡ�Irs�T]�F����≌$�%�{�D��c�UZ�0����:jƬ�ڮ2]��n�ZxtS���V��w�O���UU��\&��Z�j8��n�-�������WI莶�?�?p��B��Pu]�J9=u��4,y�k̓��0�!F��^��{���3̤7�YRs�?O'!��+�yeː+v5���BP>$��[w�v_�2��N��Q P[2��iYR��e�Оs.�.�lZƓ�)~(�׃�}�,�GP㉚�G艷����&Y8������먝X�!����K�����_�%^Ӣ�!]��ueBp��9��l��!���2-:��S09�曈�6�E�ʻM���*���=�.F ��ub��qd"~��H��[�V}q����g������02��D|�<P}*��@�-��)��� ���94.ѳJ.��ίN�9��BZ����=���ԡ��ASܺ��;���h�"�|�����L����҄x�jt��fq95��f)�}�
_א����!8�?�� �j�~J�����=)��~Fd���գE���x�V��&
�P!��k�K֫浚����2O#�}�X�%�h3���D�G$= 1��{p� ����A4�@^��M�Ss@'2V+%��H�{U�K��ǀX��}��^08�-�����w/B�G���Ќ�Q�6[���s1N�0�ז-2�s�C���1l����m�: Oo5����U��Q�����&ܞxgS��@��%�H�̅Z�x;�� �c=�|��~l�ɠ��=]%(L�!rQ�裿>w�)�	R,�3�eiӭ�2���Zl��D�8��b���f{���reDFqq�[�dw]L���h�.Zȕ1�9�}��x��Ri��1M��49L�;-�(I6�~�iC��I�-�%��Ʊ0qu�؝&��*H
54��.�a��I��#�`����!q��z���Ʋ�����R��(YWw��5xz���x�� �%G�1
�G��Ӝ#�%���N;��t�V-"_F�5�=��M��
��9�:8�����j�k��(K��y�������h-��[Q�s���c�7$��q����,��Aj�V�p��}1Ҵ��2��v��H �eI*�Z�B�'���*J�e*�x�$� � �ke��$�f)O<d'��O$�S8y����}s�I�k^�U���X�?)UA��0��jZ�:̉�=*%�VL(�z#�rk����V�'J^Ǽ]�)J4on�n���^@L�R�`D��=�pf�\G2�wN�K�L��@x���T��a���vh�^�/eưhϺ�%�L��/�*����#�KoJ��-dP��\���~��0ɾ��=r����F1ۋ� ����|�k����($F�c�~�N>������������2��ec2�%P���B;"��41�_�V��$�O;n2&9�n$�3�.���u~�t��p$�5Ş`�'qC���h�J�@<�n4{�ւg-.H�YMȽ��8N<��Z��-���^A��V�Dx���j^��u�\���rN��U�7�����]��z�G�S��'�ʣ��W� C��SZ�͋-�4��H�cI�-���y{]=���� ɯ@�X ����=��Y	�{�54��6�,���#��q�6|��%#�Xm"����
�;sc#N��pem���jɎ0so��'�ĤY�a��2Z�"A"��֤�?g˳�x�0ZO���S@�7�K�Ap��x���{pw�i�OB���T0	�,Of/k?�\[�ܨs21U��Ҵ*Y?ڕ^ ���J��?����:k|VF���y��cX�&#��
ɪ�w1���1VcLg�����O`?�Ș�q�0#�r�@���I"%��!c��D��<��=�O��OM_�IL����\��r=0�Vq�~�j�U���OYxPqv0��F�����rUf-�̡"6��(f���y���u��_�OUo,���Ϻ��F�i������,K៝��ib!�c��M�!t��G���|W��^u��jonR�:�
.c�XK���l]`+;�hIp��H��u���~��ä�`B�Y�{���Dc2�9�3 �c���i؊��E��K��AH4P�$�; ���Oӑ�Q�$��Mʟ���=�[���Rt��M��(koT��k薳h0��`�x�R�}�7\�xOl��|�ۈӵ�h�?�D�iřa�(x��[D�f	����I�Qn`>t�8����߽V�Vj�[`5�2ke;��*�>�/���v�Ļ��nfTJm+?ǫ]�J�K����v�.��d��;�M-3�!ֆ����#�C�7v�$��\����W/ZU<�J�4cM��ϫ�~���,�q�)�UeJ&�;���)w|�م����QL���&��w������8�( �	ʠ����/6��x�H>���\��(��?O���\k�����΢��p}4��� v���F��H���G윕�KD���0�+�9<:�2@U�M�1#�̏�G+��
�Y c�|�h��y���m
{ǧ��c�	?�X�v��i?;֦+`9ǵ���e�u\�����^��H6�ru�8�����%R�s7��ߦ�.�2g͗�Aw+�����{%�D�<O%9ҡ2���U�o�xkLb��4��G��p��½&�͏�O(k���t�_ڗ��E�֮}0P�����
�k�0 ����WH%�$F�qkr�ui1�}�O;\�=��X�3/���*QY�{����'!ƌ�Lj��UK*H����5w;����R����So��� x+�	tP��Ѯ�s�9�τL�y�����K��pV.�ݫ���0��V�٤s|��}q�c��8箫@/yҤ-뢽����Fp*�O��:��>�V��<��G��Z���UD�z�rĪ�  쐟�>L�P�o������w�9�\���f�z{f��6��>\��h�G��۫!�e,@+[���)��<Rɦvt7Aj:��7u�r�A��o����fQR6���^�^0��O������hA����TSxv;e '��#��5`�[8����O�I*A���j���r/���"����)�6#]��6O�^�b��k"��d@A�"�o�QM8�O)�4��0�m�����6�f9��N<'��2��W�|�U��tR��JQ��R������\��ėJ � �O�*��j� ���_�l+�s�y���;�#�mojg�U�R�9lf�+�\lF(�TFd�`����Yk���&���"�i]2K���>���\[���M���#��������Vj�#��$c��ĔO�P?=�ZL��[ u*د�S��]�
�&F�!�����arP��'Ek4G�9���Z�xm�lv�����0�L=��c����9^����&���y��p��4���ݤ�m"M����pg�i��~�\����b�5�j�(�.�y�րQ0�U4�l�U��,���#�v�� ���D�~}Qn]w+���=�������_z􆺲FI�̗�z�V2u�L�ぴ5�
(QL��԰yԇm���+l!QK	a��ߌ{�Ub[)k��i٥ag�*��o&y���a��Ӷv��+����\H�~ޅyG��ɺ��݅�V�v����Ru�BA���c�I,����?�`*���Xc�!�I�ݺ�2�lǼϧs[lƹ���/rx�̑�X�8���w�6C�lR?�PG��<��r�:w\;�o�y$*	jړv�@��@��ǽ��Dđ �']�{����ryk�=�I�^�"��E߹NȞ!����;6
�� �o�!���e{!��j5��R��#�:�]��)�XLF7�;�u�X��]����A�H���[���ݽ=?$�;���!���n6���Eb(����z�ᜎ'R��ը�% ��me��W�ͼ9�[�.={�}'��	F�* a�[��U�� �&�4���$/S��-q�_�����&UVS:�G�d�.t�k����p=
,���7���(~�6_���$K�1���D�Vx�d1�l���o�x�p�6a����t�X�{(��v��bXj�NS�Ǖu  �KӋT��Wl�+L�S���+�Y���k�~�D�����&�:Wlz<��$�&.2'���vg4�ۥ��x'YY�tC\
�/�+8�J�x�