XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������yĘ�G��a�������6`6����>�.{�'�Ҿ4ef`E��mM�vj}�`G��iT��G��
�bK�����݊h�:0�އ������`���&���+��6uȂ���g�P+ml
k���ƲG*@��L�S���a��T�g~.�pqt�O����hЮ����q ��C,d��o%��Yf���#���8�@�ܽb@�kޟHW^��4 c�����:��
�U�W7컑g��"d��_}>H4��Y���OG1�9`�����K�����0�)�0S+�(������C��S	<<���������x__��Z����XS�}ǨV�;Q�Ć%��(�x�P$�@{��)1_�dɮ��i���n�ң�0��#�F�Kkz/�z�}q�?�p��!n� ԁ0��6YY��LV����d�ܔ&O]r #���ncĭz�r�`ԋ��_�/X����B���j�n�$���^ފ�E�vp�g��\&/� r ���v^�>yW���� <)o���@@C@V�=�
���@���؛�nt����f�L�2�ۦ����1:�\b��7����)~�}�����0�oJ��X�����_j�/)���9�e��$L��HY�
o!^=�4�^�����J�{�˜n4Gt�{�6��@�M����!a�}�q6�$A& k�[0����%>J���z~2�Q�}Q!��u~�.�eP �&���	j�"�j�Qj��]}�(�˚��{4:2{$6՚EXlxVHYEB    7b69    1990�/���˄&�H�~[˨�젖�F1��O�1�@4?�N�M�� ��֪A�g{�،���A��<�q�s�}�!���ۅ}���xAT��t7󬯼Csƿ��U-}ĉ�z$Y�՝��(I�J���iU��wcl|ʾ:�[��`6237P@$��a���RT,�A\��U��؞����:# Ha�$0�$��:��h3�&`),V�=�=�19���0�l����]�0���"��
<����S���,qE�/�tl�2�-O���<�
�t��mThjQr��L��6�n�mv��ӝ��� �?f\���q��K�)Ns�AԐ�;�Gf�A�� FpkY��kY���ή���A�aϡ�T�PC�x:�1�!K�X�&<�c
�k��`c�Ѻ�Nt �[eJK�*�˭|	H�Au�s2���62j*ګCZ��85A�����ȥ%�0\��lxG�O�4 ��v��M�{J�ON24���6�t��4ya��\ޒ�e����}�������rG�U��h��
DO.+K�����U%5"V�[��%Zm�k��N�Rag�=@%ϥŀ����X�z�h�'|*��U���%�%׉�Z�_�w�b�23�ˊ��@.�s����4R�����j�$��
��"�~�7�hILs[�Jo$�q��/�ĳ |ڔ�Lx��'^�4u�x�c�?�f"�,�1�>;�"ct[� s�)�p��dHt��RD[1�SKB��z�X����Q"`��?����t�Q�3���F8+���v�]��Äu~�$���~�v"a����˱&�i� 閴!�t�`�l��GH��`�V�������ja�孯hG��:�;$6�9�nkb<	DA#�\`�\ ���ON�lXE�l6�`jO��Y�^<���<������Ŋ=9$n���W��%_ZĦ`{H��i�c�E8X�g�*W��������ْ8c�"A�Q��b(`ZD����"�������Pe=<������b�n߉�ؠ??�֚ h��<�	��W�GE�r�� �4aT1 �2i?�pj������ux��t W
�'���5��"��pZ4�p�����ukK9����,Z���)
��&Q孀T)}5��Z��:{/�n:W%[�G�!�W��J�{� ��3}��t��}F��c/��Sã�@�:��Dio4b�e܌�Pg&ݰO��5Ќ;P�R�����4p�v'��b0��V��O�¨�y�@�J�-Fb@%;��dvr�����Ƌ�P>��&2/f�%�U^u@y���GJ�f�=��e���OZ�>#DI��<uZ�\s
Y�W5I���{0Ǆ�� y'0��N;
 3Lhr���{��X��JgRS �Rj��$t,��C$K��tp�D@�Gp�q
��R$�T�9�F]�!��{Kj��0R+toG�����Z4�?��q~pj��$p��
n�ÚP�PK��k������b_�7�}͎ƦE�:�� CO��'*.��t޽��������O�1EKHX��e��
�)`�����r&#LڗT���D�uLݩuh��裨��"�c4޹��\�;Zr�HE��fVGi.��}`�H�/L?�lwk_�)�&^L����,z=��~p�q�rՆUq+�m<��+�Ml�qnc��A�[�U$d-�̌�����3�H�]͓��Y	�	dȰ8����ބy�~�L [5o���Դ�s.���OH�O��W�g���T@֐������l�fV14$)���ƶ\�#4��E�ү�+���u�z/ﮤ���~"�$Wq�Tz�(_��o�.e�Y�0�7I���B®��_�:�3|q�b��|�3�O�f�Ϭ�!gP1A6J���E�)-�*l�,�Hvʲ8�c"�\�4����6�j���>�K���^�u��� �����ՇZY�w&�}#��-�bϓ>�g[�����R�4��{Ǹ�a�vb�G����,��\�PG�.^5�V,̈�9Q��l}�&����wDI$sRQ��	Z�3�>$x�~��O�P����O���{�'�/?g�T���޸P���������W�J�fT�1���Ql�J䛑I��� �^����$Bd!]Œb^~&=V�������۴Ӻ݆(o�T�$+EBu���pǣ_8� ,M�� �����v{28r]ԿS��άP��2"
���f�TvhL�(i��l���4��N���D����NW(Ga� ��}%��OJ�(>I���]��ˤ�W�B/wLCeFn� ��k!pY�t��^�jB#��é�팧�T.zOt�`������ۥK? �#(�#�!����%o���h��}H�uV���^�s�������@m�	��e���]!�::�p��u�=�ZU戟��bE�
Y��q�)����4<d�l%o�O�ޅ$ƣ������v8��\f�<(�PbOҽ-���^t�KcO�-z�Կ'�`����"�V��&�	d����ozj�t�N���6<�-˷@Z�6,۝����輛ꅵ��������T��R��bK)�$�X��)�K$��j4{!��#A5=�������=���eo��Y��+2~7KY?h�$��R����z:qE���֡��J��mC�g=�q��@������SC�Y�j�"1��1U�)�֟�:��`/���gِ9���:�x�ZM2��O6k��s$�\c9I����`;i���	�`���s�cPv�b�M�*��u. ��������z^͠3{���9�V�B�>�]����)YC����t���;�qi��zԆv���hL(�������g���T�������72ы��)v������z25�Y����]hmB��$���J#mO՞����k�2J{D~C����8�϶�d���m0�,5��E��cs+�<h�1ʢ,{vZ٤zfM���	������167����9E�c�Z�A�D��՜N0���:����z�wz5#^ܴ���M��T�vVNI�䣭h�vB@��<
D@%���n=,HY�e�1���tG{wvP���R�_O4���Mt봀rm�������6Z:
�m����ߕ�hᩨ9�������1i�(g��@���)R��rN�]�jĂ����{&f��`������Sp�e�ˮKW�ˑ���R�ӶE��YM[����^vX�A ���|�3_@��Ҷ�Z?P�k}J
��]��;�bn�@���𺭮i>�%hP(̱�U�P�E�jQ^;&����0'���v��<�Z���P����<mn'!�%�z!�v�Rዌ�W����A�ǌ/v�ɲ4�#G	^�(��w1�8��"�xK�x�1��8y�&	����+�e{9͔�>���c��(R�c�߰�̗�]��/Db�&�`
���@�6��wèޅ�E���h���Wԡn�.�K�/v΍�]�K��ݐ}R%�pmj�O��Ӱ[��MHH����z[P��cFί�'D��:J�y4��C :�� UE�T�l��#q[��(��*uKXJ��*�ᰥ���澆fZ,A)vs�_45�� ߴ�N�8�-nʨ(�J�s���V�D:�[,��԰0S�A��Y��������l����@%L��b�4o8>v�/˕jx�I輯|�l�ʈ�׼���׎i��o�f���:����˙$�ڛj�I�6�H�V1���I��\��^e���jw3�^�d�m�=8��q�E-]['�Cz[&��Q�;r�˾`��u��aώ�u�N��&��w���/�A>/���J(�t����rb|��TX��c�[��y뵑��~��NIF�ӣ�4l�q�߆������T������i�I7ۍ��Zg�z.���5���+�6}�77?���02��7o���ڄ�X�A].k����e�,D
����m]7��(���>]Q�>����4�Ӻ�N� Zͬ�E�IL�/{��fU�H��"x��B@��g��#�5|w"����7�{T�bKj�R|FAnf�1����q�!�I.���I�r��R��*4��.��E^4$�5]1tM�{�f�ȃ�~�\ƞ��� �M'9��<��%�|ݔ�!�T���a���g�Nh��	'�FU�=�:>(��;	� �&w�8����l��N��h}���N�[�X��l�i�!vhV��cw���K9����� �������P���]�+�����/T���۲!n/�<�|���-Z�P΢�})XK�>�1�~�!;��ځ�+32���.@`V�"�J͊>p��'�"���}��\u��`���ZU2z��h�����ܟ� ������8��\c�T�^:r��8d����k��x��r�_>蟛��T���kD��M$�][�ϡ�!�
{
�]ևE �w%���P9�I�����pq~̂#�jc�Z�Z0}�GF�X���g��Љ̂����� �x�@Ri��	=_���cC./��yp�@d�߬;e�i���>L��1*]N�{)��S�6S�nXV2���|&8�z &<�D��\�9iW�w]6��/�>?�ʌ�.=�}ω���f��d�{���1(;���H�A�@���=	E~��	�.A)�ez�t�:?r��?K�ud�UBR��|�P\��g���<�������dѝ� �,�4G�p_�k��!ڈһ���%�n�D��M�0�����z<�N]��\>+=�N�
�2ģ-�+v�y�Ye4*@,����ϗ��T\�lK;SMaS���8�Qސ�� Ǚr���~��QX��#�4�����+�����y�儚�@��<�g����;5$�������%������*�C|�#bN����BI�1��`A��Ք~N�}Y����Q��	o��љ��=�㴂��ͯx���ҏq»l�W�0��i6���ݱ���Z�[q�W� �Et�^dvZC�Y��ӐÈ������Z����q�$�Ù/?�I��(I�Ȯ�]�2���7��]{����**���_t���ޑ���	1������n�����6=���RD��83}eĹ��a�>4�����X����h���Ȇ�R�*S� ��-�����Zw�o�c��]'�+��Q,���Q�����fw�%
�T����3��D�X�ꊔ��䩊%c&g�e�����6å-�v�0&ڿ�	��\8y��<}����UQ�� *&]���*��ʟs�U]��{�M��Yʎi�>����זg��xἛ=�K���̔�[��f�:�z!��viR���."V&ڐ�� J�~`Z��?�������c�<�zgp��9K�g���3�u�����*���u<�����C�V$��0�?�����W�[c^��)�G2S�0���r��~�{��V-��@�w!�)<#-�)��g_���띈{���������nn�3�:��Mݼ��t���8��li��ز�y��R�w�%�i<rR��;�����"���7����4@�e'�G3��V`�Z�����+D�a����!�z9)�w[���Z�D�$��/ѵ]2~��k��ri(l����/TQV:�(y�|��^�+���SQ�3�9�z��&�3+�p�eR��ҍ�6���2�%�����7�; u��M��s%�����_�L8m�3�_�=�G��Fq��?������_�(|T�>�S��A̼}�Ry?��H���7!(��y���$d&�ܚGA,�T(�V�J����s���D��+���"����(d�)�Ûs����_�3��3ʫe(��n�J
�qn�!܉75܉Ĉ[=P�0�?�c�W���� ����9��9Q5�I�ܾj/K'ߦ����/�D�?�Ϧ5*qŊA@J����Q7���3 S_o}^����fV������Q*C�2���w��}?%Gl2�V4�P�Y<}��c^�i�ȝ#�
�A���].8���,P��	��<�-�P�����*p�K֣�BY�>B�$�R̖�_�NL���>]�A!)[��$!��A�0���i�!~��s5�F�lR��B�qvl�~�b�������#.t��y��s�<�1ŉI���"�-�N
�q]X�����@F��2��05�M������v�|��掘3�'R���,AEwi:�	�9(▣s�c4���x%nK����m��Ma�Hz�&I�	��κ��گ�
������KK�3~W��#kK ���O����� Y����M'��P�5#ޒ�i����ѳe�Ii��'G�舔�3����1��J����/��˨�Pʆ� ���Yc�� �Ϟ�"N�LSG��" O=��-���3,�~-�
���h��W}}�b����-���m90ǭ�;��7��//'2�1[�q>iJÁ2R5� Aܭ�Mo(pz�εb������'���O�i�^�l2��yϨ�9 �Fk��'2vwX�Kw�V=�����:�A(�ѧ�A���ˇJ��:���T�\V