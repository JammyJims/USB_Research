XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P��LA8D����
bHk��!��pM����M��M�:�'�ԙ��;`�g+� ����J�x�Fl�m3���� ���|�k��K�8AQ�˴�X���,�]��/�_��MI�(�T� �͍�{�eH�Š�2e��}Q�ם&� �[�D�fA)��P�7�9\#MI����f���t�$P #R�tv�Q8�s=�˫0�LJ�1�m�Ko�]<CZ�0�j��F��.j ��^$d1N�9�R������5��av��mi��pVv��\���:�Ɂl�ڻ��Ń�y|��+V��;�N��6ڮ�b��l,4%	"����t�����w̑9��YQ8�+)�H��HU��L;�G�9�Vk.�o���S)���^kn��-i���ES�E��K�ք��#E{�H���!�q��Weև|֋?��j1� h��o T��mƅ�O��3���x�p�[>;���а;�dr�1���a��k��:����XBD�{��?9�g5p��Tpg�6ŉHMˈԮs{sc���pW�)N��:S��A��ޮ�J�P2�ɔ5�%�,���U�k)L�{3v�����#+Ɉ~@�Џ�Z�>1�8�aF0?�\Xi��F^�"g��:ŏ��y��<�\qMfd[�'�@R��XRX���g3��޹�jq^&P��&�`=�č�uWk	T��?�b'�JĎ��>���'�tX�5C7�L<=���u;�(��lp�V�����ѲCV�t�b�'��j�XlxVHYEB    4d8a     fd0n	A]�6��ƐD���|_IǪv��.a	����óH�qB1K5��n��A����Rk$b�F�mj��`ަ�u�xQ���O�w��v�(�𠊋2�LÔNÚQ��d�i���C2���[���0t"L��4�P�?Ӭ��8�����h۵��N��4�8>��c't�x��0�r�^�#��;(���,톟|�jU뫩c���b敫� �a^�Y�[�$;�� ��7گ�X!�1�}w-a�	]�ɞ�+��Aڱ��A��J�Q��>M��7�N�m>u��1��sz����*��0���'��(��KPg_�o�m�����%YY�`��KĈH����c�J , ���<T�oR ��Ƴs�Q�bt$[����г��q<�Dˉ���~#�ަ ����!�d�Q"�ն�"s�r�nٻ�k�Ry�3�u��Tg�s �D�Jׯ���<�}V��H�gN�2�)��(��a6l \��\e���u	�D���w��>Nҁ�Z+e$Ҵ�^b����7
�Ĵ��0ќ�~#��*�W����U8����^r���郘*��/x�i�O�]]�>N���9g�j28��3 ߈5�	�e����\������J��ܺ�{����n�����uJ]���x�9�{c~~��Lnl^clA�J>�)�*��=�wo=$+�;{�u�H� "�y=�R�~
���Wq���gW4z�9_�in�n�	�y��$�j��c��(Ћc����I̬ �*�E�jno<S�E:��wM����	m42��khi��x�:I��E�unݫ0ĸ�beB2MD15�"�
˔E6��Q�M+A8&Cf���� �r/lA����2NWPc���2{ �b��9���מ`ᴥ�0��/$��U� $��صq��*�&G7�!e�ڡv��#�(�~�,����a;�Џ|G��-��c�v����2dUlʆ�����3�nJ�h|wq�H�����*�k|�bo��q���ǅS�[`*؟�dkҶZB�c�[di�Ë/L�	'+ӞqS����@Lv��[X�`�����?�����{�\[�y)�wgHX6�>61��@��ҚWu	��b��w�Ir�V���j�{K��@�c%� �.a��wǘA�se
��]j>�{�\��N��=�]g�߱�Q勘#"
��H��}�/��(��&��ش�� �����:��O�D��G�d�E�P���u�M�E�Ж��zv9~��������v��3rl:�^��~�����L��֯�"�` e�t��&�sCb��e�&7I� )ࡍ�C�s�._M��"�dZ��bߏ�5��D���!,"�	S��O=ǭ�8
�3�kl�0
a����,@�o��j������$��T����dqbΠ��Q��;��K�BN�� �V�v�a�=��ҏ�0�fk ����s� ^����ME����_7)�rr��W��T�U����Z��-�/i?L�^����J�U�jpe�Bra�ׂ�5���HA�̸ZE���$�EK��K��2�՗�Yr���w�w�2�J|�l�%�?�����z-3`�!�?��/��M՞��{�FV�w9�2�>�4T��#�B6��u�~�gw��K"�}~��m�S8�P��&�^���n)C��BTƟ�F�c��2'��K���=١�C�睍+��D�qd�좆ޭm��-��7��"���� �/�e�7٩��kB����`�'����i4��v����3��&{�M���Tڮk��-�:O�H�2]��S����ꎊbm� ��j��{�#�X����Q́F������9<�I ��89�m�Y���n�����s��(�ik��A�<Kkam�ϵ��w�5�Q(\�v�:����M%7�J"-�{�(k��y&�3R�X�k�����v��P%�)V�Cल9(�|s���U�1�������][��|���h���G��˃"��B$��*�ɢBƂn�����Z�Yf._�Z�9c�Փ�hI��u����hu>���@��1Wl�G����)]h��^��'�F���G�jD� UF���Q A�R�WCGws��y�#+��[�P;��dX]oԑA�x�-��V,���'^S���E����L�+���"��y� ������n?;@>��تk�R��&嶰;\S���:N�F���S�VZJ���$�s�)��q.����l&�-���e�� y�TݗSJU��x�^���9�Nc0��QlGQ���Ik:�� �_�2�w�?I6v]���Ͼ%Oʣ!��H&�����:[��ԍ{��[.���`��i*�c4�F�{�����C��X�!�nT�{^��zt��$XC}}}Bl����A�f��6�nԚZ�T(�������'���a�g-�CA1`o
 `<���헜5��YcX@�#��`A�c��n�P	K�`6u�P��c��;a�N� 4!2�)`��Yi��V]�v�SVU,��1��u�)��.^黻�ϓ4���_��}y�zp-_K�z\��ϋ�����.������LiX�(뇝C��k��+�x����{�!�141�b�Z&=���R���Od>ٱmr]/��z��B;��$�K�Cn���qBO��f��V��[A�r;��$��}|��[I6� ,.�sY((T�[���"'���c��0�Ꝙ�5{��n_ K"q>������Kb^��+X*�QK�O���n�B�}��>��M�����M	q�}1���:?�*�݆���^����RcK�8:��}�]">�ۚ�p[6:��s
�9B{������9K���nE��c9 �Nǲ��x�9wU�:N�2Ts�s�'f���F��`S�N�9ƻ~!�+WT�ד�W�W2�)�#�=���G���l�QV�@:ʅd���.X2-]s:����3�?�4�l�ANԢK�5�齈�ZXț8��k���v�d(9mgc���C��LΛ�Lެ�5�8w�v�}��])������6�ٛ�����H�Z�#���kj�Zg���Ng=�M�+uD�Jzu����|6|��8�/>#�Pm�~s�x��>	�hs�p*�����Dv�B=Ѽ�!L׺��8Ki����������������~ݩ�Z~1n*3�/�z���r	� ��3v!�}�Sz���vyط+ٟ��#檝FB�_�hP��[�6ƴ�lEr�9͗��mN���xe��6ݫV�l�C��������ZK�{��O�2��翊�~��6_9.:'���d�\�B�M%��v:��4��i�����!�$�!�<8ʘi�����P��R��r� .q���%���#���xl���i5.D7�G�z�؃eե���ɖ�J��&'@��Z\t��X��F��������s���g1� �B#��^�5i�4��4n%��҃�>f90MR~5���3ՙW ��dI�-��)�Jh�;e��9$-XҝH�̨-�\��X�We��[:S!ܽ�k)��)-�J���Ɲ*�>b�u�L!j\D���]��J�ު�(�H�]��(�.�B�A���r|��&5�.�x�TL;�I����{�.�&F�Z{S�MA*_�m��)�aO5����WENb	�A4^�]��z��$�����D3��E�@����̥݂�$�.�D����WM�J�TnQPR%�)�/�F�I��@n��(�#�ۇi���xp�8���M�/�օ�m���}^baC&`�����F->�{W��0ܬgV�&(ߦ57Ͳ�ɲ౿"뱱��5��тܓ��@�%��4�\�Z2]�k:��(Bl�ܽ[f�� ��dZ{6AY~��A9@��$�hvl*ܳ>�S��	��y�ݙj/fJ9)����Z~���yP��z�&0�wX�Z�*U�
A֟�Y�,rv��[D�!-��lm�1�\��)��-�0�ͫ�}`.P{活�t��fac�}�[+������Ƙ�<����bi�X �b�V�"ҋ���v5l>6���m�S�"$O<g�� ?�pZ�2x