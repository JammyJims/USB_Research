XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?r�s~��?���C'��t�W	S)�����8�>D�Z��-�y�:�+0ʂF�Â!��M.S�
9oBVT����� ���]y���l��;�;�x��Bn�_-!���n_��g��!����~~��\�Y��� K�z��H��v���;ZZ�cѺƛG�+Y�Qw���O� �޲pf���L��x�7���1=0����֦�6�����?;�a��*(L/ުB!"yKđ�B�*1a�5��'��w��?+��KN����Şd�"$�i��1��{�K��[�Z8�җuߖ�$>��l�4g��l�~���~e�v��[@�8k&��P���4ԑ4/~-jp'�$ @�����%E[�F�$��h����Ǜ-�1C�k���b�>y���Cg�1�I�q��Rڴ]C�T����:ZP���BN��]��{�č�-gٴ|Y�n`�>]��T"_*ʃ��^)��T��A9�LR�����XY/?����n5D���S�#�/s�D&6,}�U�O��}�)����+NN �w�ν�����x��J���y��͒���[�}&���7�c�5��ۿt%����+�w��撷rV�c�Be2׽���&Z�"ar��f�ۡ}�~��zF�D�"�l��h�RG!dH�U��9z�����P��$=/d0
9R2��]
$�:ߣ1��>�UD;�Ay��/�@��Se��JS���!��o��&�H�8h�":�<^b�L������XlxVHYEB     a5d     340�k>��t��$���[��Vgg�:���s���El��A���J�n�[b7G%qt�]���1�3�O��<����!�|p�_�:�!�����H�xy9"SϳU��ۂi�Bŵ9�z^���u�S/!O"��>VC�>>w�[M�dR���2˂"&�T�/<���I���Њy���\K��"D���?�b�#���.��4(#�C�h�'V!�6$�!F��D�Ar
����'�4��ܑ��0s���)v�o�0���@�zH���Í&N�q����\��@�ɸ�e��x�P�y֡����(9=ΟR@����4b�J�MX��~j5c�
��
��U�Te�N��|�{(����$�\JmC��H�HkP��j���0�I8͚JEc�
ֈ�LQc�9h��j����{�S����˫�'눛�97� >^�	B��%_�s��&�+��	7O����1}:���*��U��'g�h�HB����UMj���xe�	�
��5� ��Z�FQ�_�a۟��e[?�g�?P絞9�R�N�i�|��?.�	��aod�L��F��2�ש�3ԛT��l�K@�%�-J�l[�Y�VS#��S� 4���3AO���=	�ؤ� )�A[���ʔE{Q������� 8,��jH�� �A��́�U#	a|N'�yUk��?��ė4/���_~�q��5˔j�u����N/���53~͗ rq#��)��k�mt������¹zY+����ψ�r�(�����<�{_1��~�P�K���:W���������ĳ�t�w����ͣQ��.�+�	C��:G�B�&G