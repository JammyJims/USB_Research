XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T�\�᥵�hr����LU�����0&����FR�u�=轉ic�g��IL����͒$yS�୼��{���N+��z��K@��e�Cg�w%�-���ͥ׺�Hʤ���k_d��X�x�z� �U�	�L��R����U�eq���1�����v5����=��7n4v��� +�a����(O�g~�2���ƀzg�L��g3����e����ee��|�Ɏ9ǕN�G��	TFz��U��ȹB qt!��_�A���ೊb*aݺ��.���9I�:�&=�8?���@q�h�t��u��߸��^�dnv�`�`1��Ɖ�S��*��2�m��{�K�pj��$�{e.ֺ>�#�o���<4'�(/�āݣ#j�F�7�m�;s�8��R�μ���1��K����@8��hl�Y^�����Dj��rV\TF����`��ճz椘5���oe՚�9��|wH�!����vy�e��t�M��68�������;q�_���gYz�����OU�:�;V27^��\�I�*4�I�𦫧�$`|+�㤐lM�Y�K��Q'u��텪ȧ9�+�3Śd�m�3p�t�N4.SS�J��<��u*)��Q�[��[R�[�S~�� ���K��FkK�m+yk`rK�`I��K^H�N���On���O�Z�@��+��ƽ�'���ŭ?�O����d�M�l�&�^�EE����v��u�B���(S(�~7N赻K��MiT��Z�S�3�e�p�XlxVHYEB    2d21     db0q�<s�Ӷ�it�U�j>W�d�pu,�O[�8����˨'��&�;1�.7<�<��#
�#{���9N:c�t�4�T)�A���~���9z�oq��e}{��D�I�q���B�����2ϕy�Gg��&Ra��đ�\c�iZ�s��V��Ћ	��1!�@�G:�7��59�^1����;�:�@Ho�/|3MN�񭑂������E�{���+��!��j�2�N!�W,p��HEݣ�k�E�S����1����l;ܿ�d������"�^_���������J�`��d���[��j��G�h�b)F[��:"`��#�T+�#�&�O�O���C�6J��:MW/~a��k6����}�)R��JE�|�q�oͲ?G�ҩ����3�
��-j�⟾'}�:�r���H��Ŏ#���s�v�a^�1���6����(/��3DZ�Je�11��~��b��X�PL]�d��{��7c�M���ӘE�c
?�Y�L��w�E#���e��>��=z!�NH����tp���O����m{�ŞM��r���'���4m������%��RA�{���J��@����v�í��T(�ʶoDS������~m�yf&}�}3P��ˑ��$4���z�
���U d����o�t���:y������鯩=^"!B}�[�I�s��Sz13|Qt�7�rF�ɮ],��룐W�(ތ��Ь>�HVLi���3=S���o7�oWF�	��9�+�A��|��[!��^�
�MV:���R�q�nJK��T�����H`��6��z��+�u���3��=<%��4;�[4P���#���-;!�	n�h,D�fnv�s�hb�|Q�X�Մr�U�j~��ZG�k)6)��o����n5ڴ������a^P���)���_L�js��j ����ah�ֿP�,����R5�h:#)��U��m�u�`�'��]�Rף��r}��A��`*[��Z#
��BD�����!�3�/OD����#���n����u8?��b����nGŅD9|��T:�ᜊ���9�e�*�M��=q��V&ch�Mu�9!�6{D��Aa�C�5�a�V�@����ݟ$*�*�T��/lL�6���t�s4 r�4�e���4SL}���5 �o����e
����vU�=��v��l���-e+e����펠�m��C�!@�r�<��w��B�*��ը�&c�M��e�RA��)���Ƭ�`f�2�!G	O�f�#:Gpg�\�hA	�Ҳl+q�5�Y>e��H�����X)3dL�V����F: @Zy�{2i���Y�ҾD3�#�ӢgQ~����;�ݑc�N�G�(2*T˦%��۬�m{^=�g+S��߼��]'��՜09��E%Ć��|U5��[M//o�����võ[/"B2"2Іu���s�;\{XVX���L	|�rn+ĉ{���+~��ش2�OQA�	}��;;ޛ���Ƽ���S�_�|�q�'�7�{��匿V@���qH�tt��_pa �����Ӳ'��+bqD~�WV�F�Ѵjqt�r�u��u���or#����ƄcB���f������G�ˁcCъ+�H)ĭ�yk��,�Ζ�ԏ���VA��FQBHr{�*�`<�����qk�=�%r��	�H4�1�E#��,[A3��q���0�2QV6�s�3&���Qt�S���s�UM�nI���&'"����ݣQfG�}�g�;�( i��$qEJH���\�qp�.�2�af�E}B���	1g���W� Mf�WM�e[ip>���:� ���D���P/��4�8�h��L<Zdش�s8�'{"e���=�3�$�Ԍn�2 ��7ya�ܡ���@��_j�0ʨ�3��Ҫ#�oĝ$����0y�c�-,����z}�~�+�W�х@KY݇��r���X�8̋*�7E��l�l���� ��W�/+���ct$��(o����<D�6-A	�#��NM���L"e��<n]�H}� atq�YvG�y�t�7Z���������'���X���0�<����<��L�[g&^ؒDȎ�l��%�6$핇Ǯ���
M��e�8+��t
��͵�1��d�Лycsrĥ��=�^|�L;�S�&��K��lb��p���$j;��0L���7R[(I�W�@*A޽V�F�qK���n��'8�&��yE����׈B(��x�W+ouס��""0D���ľE�2��w8u��b&A�-(�Ȟq�>���PN�DU�۲��f;T)W)�R`�����(�s�Wqa�����9Gj��.�#p���J����y�T���
�Z�ױ! T̚S��#��۲�U�Mf��t��o131�V�s���J��1m�,ws�{��z����EU�M���a���̵�`��0�h6�����7uE�ȍ��g�l�O�i��f�gk*P������qC0�����G�]��t��͢�bxc<�G�V��]0Ķ��Zք**f�u����&ū�q���zV{�f��*�^������r 7�>@�.�k��t�(-춍0X�u��>x�R�O�jDo=��@'�J����yNieoQ،(�e���+k����'�\q5�Z�A�lK�QxN�U8{|姸2�~f@���v���&�q���cE'�we��Iݟ=�P������x�0")����$m�����&:()��9oC`�Q>#o g^,S���p��7�) ��`U[>�`�Y�O��" s������=���p7�Hߗȍ�o'�k���̃�v��/�*��m���H��տ2��UƬ�0^��J�}��آ��v��WN�B>z��8�)@�8���9�0��5��>�b���j�Lh���n%���[��p���bW1	��o4��4���H1����+��{�x	��QǨ�J+_��*���h��� ��E�m�^��q`��1��~j|#����D��KE��ӯ��[L����K�,E\|��{MH258gK�hg�J���TUa�j�#�)�L��x��pF{������ ��k��F�/T��(�a���O��VPzc�Ӑ�eV�N!!��Q.�� E~��|���04�yӁ.k�Ǎ�*�Q4gh\S�m�V- ��Hcᤐ伃I2�{�c����H�4|rY�%�%675�&V_�=�SjL�%95::ٖ4o��R$�vT��&p�Z�jb�nK�m0ac��{^�hCrj7��Ĵy��E@h��}����4�A|7o&K��e��V{g�����j<��r�yEգ��4����3܂��B�}��ےZ���w���?���ƒU��G�8[VA�aIt���'v؁�>l�F ���_�X!�!�f-C������i^T��v�)��Ŗ�'T2��8$���w����up�i5��/�1��k���̡ϯ�