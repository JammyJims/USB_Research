XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3��IƌS�s7����l���5��x2L���Ȭ����/�y+7Ma�K��;7��8�ב�	7��r}�Jrs��?1���Ua�)b�ŋ���ߗ����o�K����y��̺�`�4������լb��o��J���|�����Y��&��o��Ta�6��IG��x�q��H�c�� �B��G� o��])��zq�vŜG?h�`�-]���8iD:��c���-��XU�iNJD�9�~��2�5��tOX��-N��z�v�V�/Z~�I-�V&=/�m������T� @E�.A?q�qm=���r@�����j���,h ����S��r�td$E��g�Ԥ�����L����td�s����@�@�B+������=*�J>W4�[݋EE��{|6b1�u�q(O�tˏ�Jm;
H�n�Hf5x3�6s������ݢ�dO��uK��!(xtm�PO	e_&ʥ�*Nc��B<��?�bx�d��t4����g�$һP�V��c�t��tH��;�4>oҌ�FGe�~�s�&��H����ߐ���7�K�谩��X[F4"����P+Y���õX9K��h�l&8ad�d�`e�{#����c#؛��܇��w�U�{q&�U)�X��(>G��B������G˞���冃��Lm}�=��W���Y��{�걼�5[�/�f�E�~S�`�4{����^�$]҇p�a�읔Qqx��v��(0?<A�\�"-W�v���"XlxVHYEB    7889    10d0�I���>���|����W¡�\D?��\���_�7,žZ�u��8Z3z�q�ρ����P�a��:F�� �V�j�c���%���/�^
�t�t�a�t��/%�e|C옵�p9���`�g��`Xp�?QNP�~-&��Ih:��HY��~�P@�f�mI��j6o����lz�l2ov�<�PQ���̹#u�f��p�<$U��K��kQ�����e"SI�^� �;"j1���L[��I/��t�sjȈmL�/Ϋ_T�|��Yx%F&$��������p��'vA���Z+�bR�Mw��m��=Y�.��F�I=����̞�R/$�j	iV~\�̈�N�ȣ�A ױM��׬�N ��9��üB9ҍt�|��IM�K�@m"B �������vx^�3��GhM��v�j4cf��(>���0�?���)�����
Q5�\�!hMLE��}�_pC8��S��"8r��E��,�x2�W�앢"$|P��R�3Zˡ��g'�hp����_'�ح3T�%�=�ـn���\w���->ϻ�/e��\�4A��~���J�"施�K�~��~�tJA�MTR��- �R��k��V�A�C�bO���$1������������S�Kn��DsK��m�|�\'C{I�d�,{2u[�Хc�}�x���y9����dSJ��)�f�q�ZI�	N5z/V�7���Cf���!��]XbN������> B�����N������:�L�:yP!�b>��2ښ�8C��*�B/�7��S��Bc=ݣ������I��%),Yq�f�A�i����=�Rc��"�r�M�vΆ�>�&l������|*���e��R�Lـ}�����y��g�>�|�ca�@n8%_t3j�0k2P�a$A�?�%�.r��W"mU7~j"�lGm����*�HO*�8��?�O<�T����o�h[�2�i���~��jh룋��Y�J`6u��J����{�곖[����}W�������6v���П��Q.F]2���qk��1�Aun�iݓ�}K&T=�MLW�*s֛�ـ�&�TyF�N��8�έ�Y�*8	Y@r� �c��N{?0�T�,���Ry~l�*��Ei�
Zz/&ϕ�uY�l���9is�l��y�oD��-�Q���VP�+1�8b���G��O�r��+<�,f̆�����}�(�H�ϓ��2�^W���B,!25���8;��_����H`U�ތX�*������cӤ�	�E�02��SQ�����m�f�Z�@`�u�w0�qlU1\��P=L���!F�{�ojy5R�F�;v���۷�W�v)� �� �7�G5�$m�^�A&q�|h[��"�I�z��k@<��X�Cr >,�	��ɠ�ا��FK��K��_�vZ_Qo{]�3x:Z��=���J݂�6}����/E �$.uL��c��2�4]�����U杞.#��<�'z����8_R{csaXDi�Z�6.o������0s��m��+��|�wX�+����SC�y)3df��ҝi�R���O�nU�U��O�/�Rߜ�f��A���Q�41꬛�^�p·�@���n��cxc4k����n H���]h���f��T��8\^V��x�IH~J#$��G=�,dsSYI4f��4�J�� z�S��&��4�\2�-;M]�wV��������f���V����0DۤT��K �Yhկ��vq��V�dCg�g��cz?��iZ&jYCN�\'\?��
T��1_���h�O��UJ�ʕCa�F���'r���q~f$o���lf"����\C�fy��GA6�l����#1H��׽ /��}[��^�f����{���OQ��G�ٜ�m}�$���P���2��V_��� pH��,��2���&;��O)�H�Щ��g�b� �T1�o@g�ʌK\���F�3Y���^�)ɒJ�_���4��|��7�K��"�e��,X���Rm��++��` Ț>,j \$��+����a��p1�صޛ��?L<;���IO������u�(����^��õs+�_�yJ�=ܵ��Z��gOM��H��)�;��p�g��ޗ0�4��84�޾:�!�Ϣ GI=c��H��������N�-(��Qٛ��0}�7��S5;�z��y��2�<��A7�ƪƘ4,ִ!��, -%��\��d��nw0=��IWs��!޻�(�q�J��z��g��g<���|�>�!,�NV	�u�s�\�}Z�D�#���2�v}�fv}i��u�I����HIy�_�&7��"y���m H�-b�&�I�Z�y� 2��O�����\�"]��sp�"���q�!�J�~�/$���L�R>����J!�p��m�}��o���d#���)Qf�5��(E,���C�'��J���z�nw]�ġ�E����zUZ<��j�u%�M��:/��y��Vؽ�
��I��,Ui*��r�]�8���I;GHp�'j7U�O[�Mh"כ���V�Hd-nRj���xp��i��f�Zd�ܚ���H�8�%�hO��A�a�T!q*i�ܞ��} EƆ��)����@�26��oa;��!_�Ǫ�RZՒ`��#ћ�c}��;x�����,3�����|i���s<Dp���s����(tQ��7D�V�yu]h��o�<S$Zݤk+�[q�-S�v2������E�Ns�t�&馶툐��k��fE���f}^U����jB�����p���x��: �l,Jd��0*g(Բl�a�(N��u�J�'*��-����Ry/C��襫�*.R�7��li��wM�M�ZܥrR�;�p�M��1��$-r�I���&�7�}�k�8�_EUׂ�me�7�_S=Z[s�a#�T��e��ښ�/��LX|���IN�_�㫱�)g$��"6o��Gw|��x$�gWqh.l��U�dR$�~v!��9X,T1z�u��;��zՀ���<��WA�a$P�i�Q��	 �o��eM�dyx���o G!3�u��A�(�XqI�t�2@W��Ǻj&�TGcgQ����.���]NR�;�6>1��om��|�	-��k�E��A�1�AjSo��SS��>]��ʸֆ�-��&S���⟧�ǈ̩�~6�kc:������g]�,�#;�A0�>�:oϖ��I.ඩ/�iL�f��X"c������s���	��sꛬ��\���!F�{v鱩�}FK���F��GG�O�����y��s��:H�jX:T��u���ʼ��cro�!F��Z(��}�f�� ?��mk��43��Ĝ�7��l-Ⱦ
�uUM8X���.�����[�V&P;�>��k����l��}�Y{����E�̂�@|K����(�]f����0rw{o|��~ \�&�2��X0�S��H>B�B`�Z){g3�l��Ů'��tm��@%*qR��T��ڞ���/\6��� {�L{��% ʔAC;,=�?YP�ڗ�0�e;�P \�?H��鬔Q���2�iq�uG�4�� ��#.�	�+�{l��my�����e�g�^"���.}���mj���X��9�@z�ea.`�e���@���ݪ�|�����Unl�h�����G�D��o��&N�J��oE��0BrC6}��1��@�:i.7��i�E**+ӹc)�1���p㢯,ш+9�,^A}��}�k!������EYr&>��w`���t�b��Sጥh.��s�@���w%#4nv��,u��-^�eT���W�.��k��[�Fc��I��ZI�2�͟"���ٶa�E�J�Xy�B���*�Q&K��f�"��Mg�<a�Hc���2����޺�'�CO�ς,n�{$��C��*�⦩y"��0AU4�'�9�Y\���1aF�"�Y�����4E_Ns?���+xSΉj\dH?�fn�t�{Z�0�== ��A���)ԙ��ϥG�1�U��.���2�>�������N&+z:�	������)G$m�eԞ%S�� `�f���Ab�|�ӛJ����tXvZ�$��"<�}B
��f� .h�,*�EZ~�$k<�D�?��C��tR�h���;tL�'&�v��[��O�x���-��9�Q�Y�!��GP�n/�!V����E��!�Or������O��f����[��c��u�厔7�,��r �Q�عK��ϥ%u/�ib�s:)i��T�]h�tT�W���O�V;��o4fID��