XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u$��n�a}���c��� \dY%���T��B��'"� ��a������ETK�n���yEl��[���WK�릺jK>���d��s��䓖�`c.
?9G�U#��&]��Qa�|h�R��p������t���[�;K�Ӣ,��9_�',�D�E���5�H��� ����vǞ}�rƬ�ig)"E�-�m�%WRk*X{�5&.��N��R[���-�M^s˄WO�Dm��N�]�2�Py�CQ�dr=vo�SL�{����N�C��M�̈x�ˍ��T%b��Nr]b@��S�w�x��S&��kF!��Qv͕*F^j\�KȮ��iHBL�+����1�4���0�z���g����!��bU�?a�4\�X�Bc��4"ޤ�{W���%a����(��?�R�G��)�2���"��6���o�%-�#7%&א�/f�maG�o]��-��ǻ�'&�x�>���3��=e4({я��^���:�j�T�;=>��;���,{T�r 3�iW��'� Fʪ������`�UKbS���ʟ�kl�Q>��?��
Cߪ��芨�J�VN�J ɤ�M��1�	�g5��V_�Uˢ�x-�GETx9x�����C��#g��Se��ܸx6-?�]nv�\��C	x��/ojoo��=3ȗ+��GIu"4$&����m�����ar��vt͡��µpĭ�kķV%�|����O��!D�g��R.�>�퐬92D��Z�W��l�:%��E6��\�t�b��XlxVHYEB    f559    23f0�Y<G���z�+��(�`��s2�pr,������N�BTS��yѳ����20}����E̇��V����M��K��*~�D�/�e���^0�p
ʓ����[=ؒi�GF4��\��tv��C~�2:�;Q�ܟg0Ƌ�:eZ��R�g�+"��.��$������o�Ű��r�&$��@�e��8��@L���s0n���5i�P�g�A�y�vܕB4�@"�s£��Kw2'n���r9�u�" T>�/6<�V�K�;�=븠�ou���鸿����;�Yc� � _Sg���ID1�	��Lǈ�7zy�,�M�2p'T�bE���FA�Ȑ�F9P�EeÉ����/��W���:���T(Dv,��]M�/��ܧ�/&� pzI��s`AE0�^��I���Yor�^�e-����73L��h�dN�m�r=&���Q#�f$�K�?��IV�d��;��+?G|"�c�,mY}�NN/��#���W�B�Ň��l"���ip�)�.�Al�S2d��;��r�!������cb�����+͟r`�NZ�oK�j�Ƕ5|z��l�ٳ�j���8��Mg:�~�w��25[����}e��
X4 �і4�+�yN�vɼ���sx{�|�������ɔ�:V�GpPA&d`����(fo �Q_�S�՟۩�2O�D?�"}�4�N��Ҋ���#�aE[e�x���%�$8|7�j�l#F������W\A�J�m�
L�:̸`y�Ŕ^8��fȳh��N���y�|���d�c��Cp�v�G�R�K�ch�VO��wy'�Bg��xo��{���gM�43���Jb��h��㊵S�ԃM|�JY*F^��ɴ����V�Ds���	��0v?# Z�j9U�g��&��ɂaq!-%S?�qz�/ة����QIk�BZbx�_̺�GRr��y�%w2��E��ٖ+�x�J
��;8��l�]N�p�駂)���c��}���j��i�1�ʇ(_t O>��W*�J�q��d��I���yC�R��Q�5V����]�3�|&�+��u�M�Y�����RH�7�|�c�@�*�����u��QI�y��5��{���7�g�g���}\�q ϗg���O���	܇�s���4��]Y_�|����w��lDh��\�j2z��0��p���9���K�x��
�T%F��#TU�Z�k7�2���`�ZN='���s��1x����:@��k�[��r�$�`���#���:"�e��B+K�S��R���!��{E/�=r��i��P�O:�Ѫ$Z�CG�ә�CI]�.�SéU�A2�2Gf�cr���q�����י$���mQls���u�'��&�k#%�"�z��E�n�ã��
/�o�x�3MX |�.�����~��|���j���k���ClM��HY����Ջ��
e��j��%!����XO��o3����y$�"V8�;P監Pѥ��$퐋e�������ۢ���,��0�^R���O1}r�{�&q&����u/�1�TMbOU��0�	�F���\����t�נ����_������Pn��&�=���;��<����b��������)�mz�Y���l�3gJ���S�#IŜk������I���.����&������A)�Jx"��ݮ}�@�_;�PZ�d��@S��4�^�k�^�OW�H���D�>�T�},�F1E�\�\�3z� ��Z�a�f&�Љ�X�qX�(B������L�	195�k��?s�g�a%�-�̏�+;��q�S��2%r�T�FW�5�[��n��Wt�͆���:b�H xwڴ���14?�X��~d��?�g��5�5�K2��l>;��
���>-�Ս��������o����d���LCy��i������X��0��QsC#[�x����J�����,x�6��V�A�6+68�4��-�7�ϭsl6�{c�Ɛ�I�2]�^�I�Dl4tG�)��EMp�:��|�c��"��5�����( �8=����;�Gi��|�4|+zd2Ie	Fa����<�"q��.C-E�Ud�0��R�{���ȵR���j�s�����d�<�}�uETy�
t���aw�nv��Qw�.GcӐ��?��c�#�GR&���]�b����Q��LR���.��Z���� �Yp>M�?�q!a:I��Zɜ�gP��f��D�O<e+��``G7Ⱦ~���P$Lm�|�՚�9��l�{�3F�X��*�/�YE�+l�Rw1�K����:v U�R����ݬ�N3�l,�>"%$�_7��轃����]=�HףKk*��L� ��x���T�T̗��1%1�tD�T�.���O����3����|����!���Oy�6W����߳��4{�Hȫf-��e�����c
��޲�D7#Ӧ���������YH�uM/*|E�y�Sк�Ԫ�99ǖ��)P��OQ�r���3�M��G��p1�S6L�X���h�~CW�^�
f&F��5�ex>?@���6H�UJ�W1/��}~�D!�S�_�?�+g@ۤ*��m�� uP~�Ŕs��GW0F�û������� �7|�y�<�>�{R��L�MH�+;տ�ebq�<����3����G{��Z�9, ٔy��lǦ�n#&{��L�`�{֧͑������Z���m�r,`��!�?�g��v��	d���G6��;�LK<&����P�֋4�KvTYd��:U��FK�Σ?�:�RW��3�rA!5]D{?%+Q�W<�^� �l���K6�c����aϰ-�on������*�i�gGo�"`�8���"~�`�ل˸��z?�pu%SQR �(�3�<�k�O�������W���p�YmNL��ȩ�d��a�����y�׃�U\qS� �H�U�=�e�����@��M&����XQ�'eI5� �W:5����w����[������ֵ���Nf�OGӣ��+���du�mx��+y��}�w%N��3�6�.���JX������m�=�\ ��� ��1��M�(�yt*~7��g�Jq9.����J0�l��������%�s-;��t��~�]�5I��v��@E>>��ݳ>E,n�Y(D�C`���W�C<���cQ�u$N.��R�9����r��h����}*��F�4n4�i�|��&���ݮ����,&�[Y-XU�"�;���n��l�&�*U�(f�$�y�y�=Q���ͮq��mMT￝�~τF����޲����0zї���7��ׄ��������&	P|����R_z����,��r��+y���T�:��tR���lv����aw�C39����&��q߻A'E�~t����5�wE���7���k���r7� YX~k,U�KS�V�V�^��	~��8z�%����2�dW|R��D�Bؒt�$�Yk����@����GK{��u��"�2�mp4�	r�q�_�V�>+��4}6,tԬv��K}.ŏk0�xE�?8Baa�3��/��y�(��R^�<�$�*]m��o��(p�� A��ek�/�@���G�oJ�.`� |����v�"H�N�d�,|䔁s%Q?k	Q�5�Zզ���J�/�.V�q3oa�ӽM)�b
����$#�R�m��w޻�	?�u&3��HY U�QP.����F~�0V��N�9�|���+e�u�O|�K+���h#�v���+ߊ��/j�R,���Ȏ�O��,���PO��Fr%᩸I��n�>�k1�Ȫ3��r�F�څObU����q>2mF/bVK����cÇw��bu����O$���ɊߧŐͻ�����"��7H��ᶄы�J�kAzL7�����p{RУO�3�
JǷ�@f1�;�wG� �<F���R���e'J�ן,5�|�;�Q�4�2���H������"���$���^��Q-[�, �vR����K+⚮�O�B�3���/��{D���4���;ˈ��JN��QG����DTy�ϙ��)����6����\�uv�>�Ts.ep"����?�!�$p.o/O�;
�g��o(mq`&���$�d��X��}p��z��b]���{ؑ��&Ķ16����Kf��}����P�-4Vb�':WD��e��4��;3~ʔ�
bW;���W����
|K+�Bu����.s��I�3�|�HM���0�H+A�3u*$.�^�`v������y�l��z�I�Ӊ��M_wuz�ں]VR$��L]����4~{�r6�Y�k�Z�{�:�]�خ��`u�,���A�#ոrH&�4��b�w��=�4s���?�u��:�p08��Z<���  ��6Ǡ8�ѕA��x�t�e�blޣ�zߴ͡D>~/�#]튂�%UѪ��S�w�V��n�켼����i����ZS�,��t�+�7U���Mr�9�C��F�l�hI�����@>b"*t��8�!錵��cZ�a7X� H���9G�6F�*:#%薬:��;��s ��^�����)���'8��/34Tr= :a;�t;�V���m��xD� ���cmc�|,���.h�Y\Kj���K�ra���	'���)�8dP3��pT�m$(���4�#ZZh�j挻?��E�b������+�U���+lap�i��5ӮdЕ��5�{���A�m_�H~{�[���q��yx��j�gҁΞ�Pӵ�����܁�v��߱J�<���K��0�+ct#�so�4�?���c�]��唅���Ȗ  U��T��AmU�CtrBi��iVH����yo����`�=6�iC�����?/v����)�Yh.f=	�B�(�����i+PS^�����Y����8����ݧ��</��O��;i�+S�Ev
B�+�n�m/q������R��5�B�B�d��8���*��Go5d'w���4ʵ�R��R֕��ݰ�B�N(+�!A�`�$�ޘ�}�6�"'l�&�$�i20֪�N]�1Q��z���]���������,t��
6@i�ߩ)�y��U�=�'�=m��G���gR8(?�\a��B�Ǒ����$9���BXpd�+A$}�fK�D�j3�H�<����dZ���7t�\�nB���!.�,.'��<�*�y�?�|i��I߁�i�=�:���4|�����Ce@q+b:0.����p�����`�	�K��bh�U��E��wzK=)����e֐u�������U�f��rv���i�J�b2F���ml��m�A�Q~�TX+���W�߽���>�[$�nwna-tݾ|y��"��������i�"�[�x�vrF^`�)�
��;��'��f����Yԍ��c`�]mq9��G�����b"h2ް�.Ѥ90�3��.$ޫ�ny`cr�j5A�L
�$հ>��dc�V�ޟX���c�麊��\Xo�>Ig܎.��ܿ�'�)^m/D���j��%�أH��|~Õ!|�,���Ql�d'�`h���Hw�3Ƚ%�|lEKǽ�vä�Y��)����DY���bz��%���砯��Y�߭E�4q�霪3v=����YY�Vj:ԛd��c�����
1��!�Y��n�P��Mp�NMyr}OP�y�����9���&��'�d���bͮwQ�����eQLv,���M=e����S��h�օ�% ҍ
 1�t�{JY�+c���iJ�0c�:n�E)�3w���a�B=�!�����X-�C�	�)�]�W����1Y��2\�Y{��5��������-ѫ�`aCo���[��ɗH�U�n�0Q<�ˤ
9�O_�
�r�����>䉥�N��R�@������6�K�܀f5_�Y�:��fo��t\0�E�Eܖ
0I�RS2�ҫ�����K-ių ��͚F��"z	���a>s�\<��ݪ5���V��<Qp�8y�?\5��X�?PzDQ�%��H)|�J�Nl5�`KMy�Q$���x���F���OBB����-j����1��q��4A�r�%	�
��U�T���g-LК����KO��4�ha�J}|��@�;D�)��V�KjEL��V�ڙO�殮����	vj�ۂ���C��Z��{�;�]����G�r��򲶸Y���n��{�,�uӥ��X��s���Y/�pN-7�6����(��Y;�Z�,&�����q��]�'� ��{�
��8��/��6�����F�\j�/Pv�ԨJV$����LD��QfЗ�QO�w� �T��ѷߒM�g1#�e,��F��zC�R�6��p�X5�	ad7jn��F����Uo�pE*��BWۺi/��Q�׶g�z3潵��g�����*�E6Wvr���# �a����khP�r���!���N4�``u"ףG(�y&�����&�%>(3��	J�-d?m7sӾ��?D�����nl�w��2�sۖ�:h�#E���Ҽ����g�&��(<�ӎA(p!a���(&|%�Kc��.7�(�.����P�\�|�s��:[<�;_0��9�澪@�%�hމ����6��9�`sT.ðHf��ʫj�;|����O�q�bV��i ���8(ݡ)�hN�6+o~�U����)�޺�)��I��`r������݅�����ov.��w����� ��;:��hV�y�s�%�7WF��"����nZ����&*;�j�in���z�SF ?}kC��=i��[k��W��hE�i��]E�-�{��\1o���#��>	`]n̠�w������7Jl'\s:���[��r� ��Ti��h�M�����ڋϋY�󑻤J��g�����X'����&�t�09f�ED��>����|�9��f�A�qu+9x}�X0�L�q�,��hk4�Q��(uG�R5?���cj��"c�5"Fi��gs�t`d�C�����˄���� �ot Ё'�9�X�����.D1!I��$HD��m��w�;���|9%2/�Z��|Nz�J����	�+�%�?����hN��>o�b`ٍ0=��>�40�-W�7l�<)�1���4f�U�#�]:5�`�[���	:Q�C�- ��x����}��>^�a#�����dz+dC����_g���	��(Ha(�sO=�EnB��_]n�`���N�i�1^�������9˨@�0?�c�sp�w����*�F�x"�E]#�9���;%���5hm ���Oy8����Ō����ҍ>���$�\$���&o}8ʕ9}�7�&?���a��.���u(��b��0 ��H����\���Z���pg��m�@���*M�V�t5BY�<�O(ao�(�m��-��%IjD!���4<`o��9�UV!�Z� ^���'���~"ͯn����Ό��ͧ8#�0J��ou6Q��g��)<cz;�R�"� ��Y����T ���^�𨒌��)_&TV͊=n�Λ�-�+(O0�q���E����^f��Ǉ�����/���~��9��K��:�	�����؇5]�(�7"v�#�h]�Ӝ�i��`�,�=A�.aXK�7{����K-��F�ţȅ^6e�[]9������y��ؾ�ts*\u���S�$��dyM\�B4������~A�p_7�_r>�	��aH���9�~)�hx�B	�0Ց��H`�p��r��-,N�=��b��R�����M�(=|�g}�VK���t�l�}6a��,�������u����tM�v�^�ɬ�&ڼə��ݽ��5Q˷�
�YJ���X"���
�h��cX��V�N����}@����Aڙ&e��vL�;��_�;U�%w�pG|#L!|��i����97��<lm܄��#�F����Z�g��D����y�^���l���j��f3V'm�t�C\Mne��A'!(�*�p=mM>OT��`^��w�2vU�D]@n�2ii5����h��|�)�������4F]T��o�<�r�dr>F��`�S9��$�-�!�S��_���U�'�7�	F�N�EC#.q&�.c��) �r�����_B���޺�l;��!U�[p�X�V�%~�U,��{Ȋ(�C8S�Ó�2�e$w^Di_S<��,˯b0�'���B/�@t�׌r�G�AYҼ7#�4;벫o��6R�~�Ǧ��K!������;���%ݚ��fs�M����mY�a��t	5b6�TD4�Z"w�F��JX|\�Qz�#�̵6��e�a�� �$��% ���W~�.3�'���H��TӹnNw�t>���$�Tyi�������S~�Ŭ���F.wq<
�jR]T
�E�("�[ӟ��̈�dP@N�2�5�\I�3�yf�Y�V�3�����x&��hu��,i<~�6�����$��HOJ=<I �O����.�NW5+lm)iyڤV�������)��j�~8���݌��~j�^`�4\p�W�G�j�4���Dn�C������G*�' ^qm�	+�.�M=(v�'*o��k�*�r03���J�Hc1��JwoSJ��J�_�i��g@]�҂�,�e�H�0!��xw����t��	ES��"D�cA�;�x�]�P����u/Az-Y�r��4��J=�&�~��g�ȍ�yo�Y�>KHB�A��/�� �}y^��r�KT�N|�_)�C�t���u�IM�;)؋��ƙ��+y&���g&W��q!|2vN)GM��s��<���,X�	/7��Vs�Ƨ�}��B	Uqzk(.)u�2�o�)絡�ȏ��|����?T����,�`����M����<D'A�L��]��8�� ��ǊiLJ�N =ڻN�hp��o�90�"���V��c>��{�V�x�h�N�sA���Иԁ��͂u�nFKRP`�+)]���ا�����e�R���.�)(�*���P�-�@�W��g�����E��&Ixu\9�R���=m�Mn6Y?��q'� 2�P��g�۴M��u7>]�M6��]pu��Ij9�$�y� �8_lI{������N��AT�gk�j��(�s�g��m3.�z��?��7�E77��a$��PBUYs�~��?t]���E�6E-�