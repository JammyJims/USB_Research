XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z�j�lFc59}DM� ���3zp�o_���6I>:�)ۈ�7H`e�nVl��(,��A}K=�yJ���I[���:�1vDn��$ӟ��(�M�Is�o�8rI�eY?Dh$�/�4_/˘s�;�@� 2锘�!�S����_���ۄ���?Al%I9����w�-��><4<�Vo�xv.���ّ3�;�Y�;, x:����﵂OJ�-��ݣ�9c�/#�z;H���;P=�Xo]�j���f�v�������d�pA��*�ڡ�_����qG��p��]:<vR�F��b0X�b
���r{��P�ٞ���O0�<w���8�384 넼*��F�r%yP؆L"����Nk�
[q�r��qY���ȸOڀR*�@�M�/��%����Ǣ��
���u��w�<*{sg���Ң��Il����Ț��/#+=�^�k���\(�2.ۄ�����.
��������#��K_��]@�� ������&��rE�H)�{k׃�%�9V��-,��R��T���}iA(n�&�))�K����.�(���J��ݶbAJ�v�j�^_��k��%blS�w���6u�����q�I޸�����7J��"����8Ꮩݑ������/%OA����	\� �w�F��']�*P�e���H��N�L�0q��:x�~S�d_�1)�?��8��5�
F���E�ҽ�G,qmh��,�=2a]>�L�#��0�@�n��,�`���a�JXlxVHYEB    15d2     830.d7�����}2B�����?���2����v����s۠rh���&D�̠%,���NM��'�Rt��bH�J8p����5x����)/�|�{T�|N�KV��*܁������Ac�_^ڽ(�B�TÈԁ]�}�	z|��������8�*�nӔ6B���6vn��ݣ�x	�":��OE��0�m����~�
{�<�b�Z�r3��F�cw�-�����*�Fߊ����:�v�\�r�
]� ���,1pP�Mԭ�-O��'�b��Rã}�1�g��p��ha�4/�m�\�O����n7�e�Hy��<�a�/��o"�1;��+�*H��
8�L��H��#��s
����]�l@�΂L;�j�T	ɈI�	2�2w?�-u�6V<�����o
����&�pCi�3CR ���ʿa���5�@Q�6���,���s��=x,t���h<��w�H��|��M���|�@)��A�8MY�p�K E�`e/Q�z�,Z��P�_aa�~+�^C�fݱ���1�f�b`Ē�u�֝LZ�Y�~��(�KZh��T����p��sa$Q�"�M軵~m?N�\�Mt��W�W�TL�鼍�͔�nI�;#1��\_������D��Ҁ�`�}K��������
q��� �#KNsX���_�ǧێ�pV)Q�ĵy�|��3��+��N_1qOY��,��x���" Z�'4c��&S���I8�jX��	�X����5L�[�DMM�;|����;f�T�󔤊��t������M��G8�w��e^s�3�9����ϨTYc�����ٱʏ��,�ŰO��bY��Aݰbp)��s'�e$l����D�Ĳ+�q�|���T��i����>�Z��0(@D����3V�u	ú���Z�"�H������"Id$*���9�؟��TA��&nr�P�q[�%8�F��K	�-�kvvYvE��� ��� ���0� ���0����h
rbs"��ik�3Ro	�^^�c�N
U��O���NdFIi��Ʌ��Sp�U�4"Q��L<�n>�;��`�iAD��)�Gr� �9h�F,8s����v-f��>b��Z�{ՊLI$\W]�R�������i�����??�JMI�
V޷�{�$�%0�Q�I��Uq*&{R�}0�����b���m-���@�3�F6����Qr )�jȖB�rN�uu�UP�}�������{S���X�?�~#0���rc���<��!�S�S���j#�l ,� �+�B<+Fx�O�����ҹL�}q�+i��Ϊi��� !��m7���8Fr�7)�^�c���_wv����C�Z`ɩ� Q�'-�-4�w߽������[��i�+N�B�K�,�R�~�y���ll�+x ��7N#.p87xv�Y����U5������-�%���*S���Q����؁�ev5��u�!�=Ő��`0�w4۲N���n]��G�B���D�� �*�g��͡�,ppD�+��]z9� 6�VA�\�1�wa�upfq��iZjN���Vy.��0�
�(�ja���j�뎱�_����
�I����T�_�pB�&�:�'�1ǱtJ?��)ћ俼�њ������"��l�X�e�'Qm�i!��';Eh��Oq¾dq,㒔�����ϔn�6&��[9��\���6����\�}������s`˿�獥����vӥ�p	G'��^���W�[�|/�n��;~�buGI��-���>��(����Ā�^VU���@+��J[t��p� ��#�% ?ٞk�U2y��3EW_iI�*������v�+�FӇ�k�`n�)��T��A���>9�J��|�+�~��Jp�(�Y�p'�J�O��Gخ�&����ҧ�;�"�&����Uy|�����xepq�$S��E1��H&d���0\�=o�R�[�0�����	�P�Fk�~�\ۉ'\�0"<;����y{0�sQ}���~ ����=�/v���S���A��y�&`�/pb�)����ͤ]g5��T��<��u��-���[-�O��՜��=/4mB��`�x