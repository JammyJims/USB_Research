XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���_BnxrN�W�-�B�YZ�����Z*p:Z��$,{��q]@)��^��jE�&���)3��x�|��n7+:��8(��hx�1��N��� �V�!f%�����E�~�绻p
Q�}�H"g���A�(:����L��	/�DdhU�K�rH�o�EЇݜ�ڤp��I	E��t`�<'8������^�!|ވz���RY�/s4�\�5�y}.9�|k�L�ZĖ[UV{v�6Wg�|S_���J�c�ȶ,��+�{m�[�+�,����
4	dzGww��$msD!/H��D� ���tӌ���֐=���w.��Z���9�@�hUc<�kO�3 �^Fu�*��S�B��3&fJ���d�	_-7&��_�`:mNh|Oli#�����r���o��D�D@^�L�Ɛ���Ʃ4ak+�@�Un��Ů��$+�������:t�O�R-���p�q�w���țR�4�7�ɂŎ�'C2�����UN��� `���A���!ܹ�fL6���8�L��XJ�yVH�84|�}�䣳��ۋs"i9ӑ(O-�o@�s���@Y�֊^{W��� �:�.�TVZ$�s�lZN=������&�%I����N����]ϑ�SST{��Ŧu�J]!"q�PW���AzQY�S��Yd+/����[8�R�V��w~vM����ǬŜ���BS㐽 $;3��'2����4�Z9��𳆖7x��HQ�#�9�e�1��+%ʬ`r�Zz�&�aou�XlxVHYEB    fa00    2940MGT��к ���K�J�}�o���`�!��F�7^66q,�����8���`4�(�=��ǸGt�����Լ�CM�h�%�o.1ǅ !���qΨQ��/��S��(���"�km�/,<���ǩ���|�W�/=�0&�� ?a�f���VS}[aid�l�����ͤ���3T�Z� ��'RaڂNDjjD>��7�u�΁�*�+���F�1dg8�J�AŰe�c������.Cq���X��|?��a�}]~�/�:g����v�)�/z�F�
6�@e�3>a�%�mg-
�g������T==V�?5�=Ke]r"�"E�56s�����Y��jd� �0�����'&���Wp�Ҟ��u��x����Y�8���ݟ��l��3힢���u�t���i���	'�cۀ��>Y$h�D�0aH��d0��#��ir�dqĂ�������6��
_ )r��,��5p*����_�<ۡ?��q)�	�m���-�?��R�$uǫp�z��Ǔ!�J�Z�x��?'5��he1��c�c�����E��Ou����x/�m�4{�Y��H*}��Gxo)��
�eݽ�y�e�5�uT�)=�s����E.���Y�K���6�` ".��K�I�9�zcN����PNջ��.�}��
ᆫ�VW�L��6p�s�UG�|vg*�i3~:�a�V�NRzr�������^=7���"*&��Bǂ����<��b���nm����
� ���.d�}!B�r�����N�i�a'ٍ�Lj�`*<��bN�B��PP!	*&��mNϚy�稲�����_$�����@��?%ϰ�w��ҫ�
�Aa��e=�lwRSZZC�x���A..�wG���n�f�^OR��R,�w7萼�V$c5`��#�B�����oՙR� �Ғ��I׉F�Vh=��Q8�ORx�E^\�l%�#�*�+p)Z�5���k�PJȫ,2��m�	�����F�e���~�-.Є���l����Tq���o����0�S>�(��4�6�8�/����E�����j���>�@�LU6l߬c�{���\���;����\�c����)�wOxhe�e�?��i�ᕗQ<�g�jt�T�9-�Y�2g�W�YȪΨ(9)|'&�8��ԫ(�����':0�r�ڧ1*$��$6��e5����,��9���^����Ty�s�����Űԝ�ld�/��$�#��ϲIG�`�_ƌ�a�n�7����C�y��c�K����8��U?��`���1H K�����EEYz:���%�czO:�Wg �w�[�N�
���|�������ö�7�/#����\2l��Ik��`l<=:���u�$[ج��q���X��za��)��Cv��&�~�d��sXp}bQ�x}ݸ�GK:��%��SS{t8
��U���K|��1@��|u��:%>�-�R�#�&��j��ζW�����O���ǅ���o���!|tuG]�s������|]�Q�m��\DU��&u�����#�4ܑ=;cj�#��hӹ��F�+��l��W���q)S�2��~�|t�D�DR'��d1�ɏ����C��pgߪC���(X��b��ӱ\��f*�&�a%g�>t��7lq�
f��k=��X�@IP��Z�(�n}��B}^-ۺ����Z���ʨ�DY��U�D0�{�={��'{4{�w����ml|)��]�=�����a��ٺ�Y���s�������5A��F�\����Z�P�"z�L���A��,
�6��%�C-��.P8��1|,$!��g1ȥh� a�9Y[~C�`�����q�<H�bgˍ�$Bk�L��V��R�m�"h��p�@�i,�~�F�e��Jm�������ם�
��z��lz���*n[���F� *}#��s��2�\����)\����I[6[6���� �_W�6�^��?9"G��T��`��=o_3�4ٿ>���� EѾ�g�~�HUd<��9񝕕Ep/.:0=n�<�jP��O�wn���ȱ%\�s�ќ
2d��Nǵ�`��_��>8�b���<���e�:\��]n�?�1h@�8��� ��pgcw���_d)��X�J�b���L�#�/T�m��>s�)FS������9�V�J��-/����t�;^F�\�ӷP��Twaf�E�6n���2�2#� ��1��ʷ�� `�CKmTޥ�lc���	�Zu.���t��©"�A����R-c��!�CF�S���LaJ�2|'���ͫ�?eu�%���EK�Ӗ�U�k�s�z=ڦÄɑĎ��@�d��ܤ����W� B-��m�,5��J�]d�6<���(5E�x�yM�b	����I?RY��]b�w�I�:r�-�M�yp��۝���
���r�E�KUKfØ�2�u)@�|�w3/�Z�،����){����Rk�4��>�k됣�*��ל
 o�]�nZ��&8��o����f
���ukZ��~@(U��Њ~�M��D�uNY; L�"�,�A���CnȢ	�9���:Or!�{���eWI<̈́Ye*xiuGʓ^k�|�%~-�y�y��Z�5����H�r����\r��v����Ҡ� 0���C�h�ޣ�@q"�u�eXk&'>>h�,���}����H�(b�D��oPP�g�ZK�ϡ�����.��F �Y�.��[�U���֭"D�pM��2=YL�P�0�R���\i��Ԅz�MD���&���ɒ ��xHߴ��7B~���3�f&t�5}�.gŚb����b��=�D��+B�N����)�I
;�IK[�`^~�&�մ��f�Y��-/�Y}*˩�5_Ԋ�r�* h�ms���`괢{���~E+=���$<�撤22�E���K��u��V�j:���n���u��O��]�
]|���K_���0q>��K�t�����p 0���&<C}5P�^ɩJ��I���,�H��MH�C���!A`(֯R'��E�������_�˅n�Ny�)5�J^g�ZBa�J
|��MW����2&uM��?]r8l�c!㖏ܸd; 'A��X�=����vsgq�a*fX���u����uL�Y�)�'���*���9��=2�-�r�=z�^Ħ���A�Y�;�#T�U��抽�V:O`w�ۏq�X��=Ă�0l;�H�~�~BC��Ő
c\������ἢ��h��U/*�R[���؇,���u4&�K
VW�u}L��1��̲��Kq��0zܢ�B�1�Ă*�%�y��|e�"���56)�_�=�1�0Ƃ�������Qڜ�'���ˏ��R��ж��1}��k$@��Ô�	�1G�*��-@y܂uBT)�l�Eτ�����7K��+��"�͜<i�x��I�9�{ޱ�i��ͽ��mb�
�2���
��'j:�� ��Z��\��:�0�^��2_�ժ;���#�}��Ʉv� �s����>��v���5�J=٩��Z?�~��*o�]0�°�R���#-A�?p��A�I�4�u��H��� �[X5��TNK�E$��opc���p�!��ga���K%1'4M$I����2\�!������R��(zѳá�o�&1��z���4;�t q#����	5N{y����Ult`騷����V�޷3����'�|lzN^��mZ�_�����;��L1����G��v[�,�ۋߓ�kT2�~�bB;��57Px��
��(}J���5�_�+ٮ�YH6���os��FM��)�{	ZЌz�k����ly%grK&�_�m��z�Oj�c��T��d �$K2W���1�@ �n�"M� )'l	qS5���uCX;|�yb���T#��?��X�y� �4��%4�g�����|�1��>�ʥ|�0�	N)c��{}��[�)�hi [�}�J�:4���2�
$������9�p�=��G�ƹ��R#��+���<�-a�X�/��{6H<�m����u�$������Q4��g�ľ�5���{�R��v�]��9K�����hٝ�K�NL:R��X�LŞ�}�.{T����Kf�$`[�LI�eRE��h-6Pȩ���/^��\d9[��|(w�7�A��N�C���u�ɴR`)���("��X�Z�FTf
�
�͎�r[������GY��28��;�y�!p�Yv �Hy3�����ZIt�'�W�m/��I$��9Z\�l�e�ތt�����*�6b���Q���k��� ��J�;��0=>�%���D��V�i��(r�: bI39��I�$�XȦ7��q�Cth��H�����U�>�,��#�������֑�gf���잊n��ϔ��)C�(�ݜ��X�f?>���6�ta����V
��u�ž=��[�P�B��\Kf���~T�T�� �و�z:���r�a����J����$p��p�j��|^���G1�*���?��7�xv	���~�?MQέ�m�~�$�J8z���J��-����e]���lx��
�o�w�[k\*lyp&�@���[}j���<E��!����yrqN���GZ{\��\[�ʓA�a1G�9��׮��ܖ��Z�m~H����vl��X.�|�VT+��v�m^�z�X�p
��4���&�Y�T�]�݆lWE]�6Z���F��q��D��P=j�í=��,���x@�&ğL,><M���>t����p�w=����i\���l
��|*��@�)�C���z�����ivX��Z����rGT�Z�'��<�=N���G��[?�^@e}��2�������+q�p��W�.�f���/��� !eާ��u#:��C��Y�� �Y �۝Po�b�'��}u�v�w
���)���;<~����
M,Fs��:ie��u������s�+�)���N�����轪z\���xGR��e�B��A�񥑲��g��-y@9�����?��W�C��I	����*��˄
�vMr�9O�����I��m~Y��1�-!��o�ߞ]��ec�O�W�^)F��?�!W¿�W�"ɭ�9Ζ`Geh�{ޕ�)��ep_��^�Xh>��Gv�s��%�Ż6ru�!b���眸� R�zA[����;�N+�;GSL���~e�<4G�^�4��8���6�y��,Dq_!#2�-G��<4���X�/���<�+�h�~`�����X>_�~NF���܀fx歾�0k'	>��^�s*�a�bG*���v�H<�J��O�H�[m��I@�ZIAP#�G���r2��í����#7|뇉P���h����F����!���m���)_��~��d��h�V�m�0��V�@R�h}���(�kʭ�1�����[�]ך��s�.b�g��<zU�dw����V7��i���M�4ّa���ď� Oc��݀���ñ(��b$q��F����׾VR#g��4T��0 /�t]�f���ۂ�ct��q`���s��߱��ɍ��)>8�.��"�'����=��L��)�u$�nm���-<��󎎼!�(i	"��`�a���d'�k}�I���|� A5r��9�0'�s� 4b��*M��dm�)�pvr�¼�:q����Pp�B(�abc:�R�a��-�bM	1�o'
{4_[N�9��FᡫC!�n�d��2��ۧ�6�����g��E��^��=L�܍�.RTH��!�bw.���K�2^
��t�jA����.ܓXGT��w�������<�t!Go�$��m
	`I���x���!�\��f�"��-�C�e��>x[Pg阀|�]�:�QG��!�i�eN;��"~�eB\��"�\�5�'�S��]��uu����x���((H�ѾD ?���қNG�R�ϥ Č���Y���-�
r[rV&�t-���a�̝��cF�'�f�!0h%�"��M���xwIA�_�%���+?�)\T�jN׫�	�{���v����9N�۫�T�i(��>��J�6��Q1p��'ܿ�~�BP/��V���[I�� MPn�v��lB����C�\�!@�e��ӰX槍7g�~�B�J�Da�6(sQg<\�p�-���R!�<�*g�E���uⲘ�'���e����25��{Zv����j�>Q]�{�l���S�\��0�C�1������b�smQ��g��k�^'yIu����S�i����ЫY�f�M;õk�M�����u{�\׷��xp�O�y^�,�ㄖ
��QVcEue����
������}��5<���k^TC"J�um���+��2Y����ǇƋ��BM��Ӷ*Ԁ�)>ƚ_IL{1̬)�T���X�7_tJ�z�$Zx��p�i���ȣ����:�lbN��))h�I�F�y!z�-�&Lk"G���-({-9���i�b�N��]ߒ$�*	w%Q�%��M�YzN�-ʬ|;���9�DWCa����m���<%�BX�;��n3��8S��Q��Ó˃�������[QX+WWZ��x&�ٱ��O��,� �T2э�o��9{�sQ�>��`	�*g��e���h�f|�n9�$/r�Pb:�ӃV��a3�����9qmj�E�K�u��i`T}��Ck�=�צᰅ�JP�:�qSfK �� ;?��cT�ǧI�Π��i4�_c3�:
� �%|G;��@q�Eg���⤅��3�̺�ք$c��DppwN>�#���{�S>����7����h���ŏ������,{�8?�ۺ��.P�0�,�����+37�U���(E|��3�7>I�5�v�v���i^Byc�M�������������O(D�� �@��7k�(�Kj�0�J8L�)>�+{||r����E��5ޙ�hS��1B�x1E�/��-/8��IJ*������u�1�B��ˌ&�6����ѪI}���A�Qo��EFU�6j�`\e q@f�A�	_�+�� V������/[����&#����jZ�K=�E	˗y2�や�MN��.�=�v�^��	��oh����p뒚+���h7pM,�d���\�db���H�:�۴>�%1�^����ņ���ݼ���k|4+<����q����a�n�nĸ��&��+�	���*h���8�x{�
�A�i�0�8�9²�⪅��s�{d���Ϊ�O� f^a���n���2�R�@� '�褲ߧE"q��Y=���m;�4�1KH�cGP@�qT� Z�[RC)���cL�F�:��岸Ш�0k�B.�P+P��A��^�%�҇�y�_eRK�]��"��t������Y{����}D�����F��	%���}�H]�2��|�@�ٍ��;��o���p�D������6t_��K���At�a�fM��+r~�ɞ{�2e@��b3A��Ւ�u�$
h$��ƨQ�Zz Y[���&j]V�mC���)cޕ����-̚����d[w)���۸��-�.�QL�RJj|���J@���R�&T�Ѕ����r�h�k�l��
�7�EkC2K����'��s��j���G���ݘ\�]��94�<�,���.�k�A��e:���*�_���=Z��P�*�lVӱ���05���4�����A�2><���YP�C�!X�<��e��|Q��٪]c��^h_L9�f�9��fu���0�˛����&��=J�-{�ǔ��s5q�c��\gGHQ���G�݌��<�a��y}���	����>m���@����h�A3�W� �9��x�	�Ij.}J�nsa��4ˇ#�Yz�z����ᾩt���3���6�M��\f�������]0K�-P�� qռbc�,�8O�LpT����e�r����Y�S��73�?-0'y�%V�+��x��@�1�@� ��|�A�����:����;a���a�R��sd;(��Y+D
�����R(3mOP-���3�!�(ٿ��22#$b<�r�Lw�ā�ԋC��ݮmjٺ[�g�E��)��ƀ<5o4�iAg��
8�>S	ú�Gy����h��������7!8�Ħ��FSO�>����/�F��Q4
�Ļ����b����|�2��bh�HP�I��)���ÈT\Aw:B����?a��m8X!�e��BP>������e&T���IB\�t�4�=���Ri�6�>0Bo�M��g�ˏ�Jg�Ǧ'��ˠ�*h�{�	���i��#�`�x!/p��݇���Ip����ݑ���H�)u2�b��o���#��0�x���H�+b�W���"Y��ׅ�#R���HB��8&�k䜟Y��
��؟����E�����xl2��O�m\�oi�Ɋ�����7�g���b���ch���-��{\0���{�{��7�4�C�Ծ���]H�� 5	� �"��X�ex#x���?��M|����G�߻��/1���ǘ�vU(\
����\������gw@�۽�9h�KZf�?د�6�щ�����d0���e
��ʰ�)qA�21vo�L����+�b��\-W�*!Tq��#*v��	h9�?��,�R(�rc�b��`�v����'��0N�M�L�'���,Li�'\5q��28���5:2��o�7L�/��k���M߱y��_.
cy.9����E��n~�^�U!�����ue˘}������d��*s4�m�3�Wх�g�ԠE��˧z��(�[��ǔ������x��i�k�M��Ӄ>Keq��M�-��N7H�ȷ>2mZ0ꥱt��J�`�;�b�C̰��<�J�����,�����6A���qW`�6
��9�}�`I6x�+A��"�\��'�J��!D�\��1b�$�:�{�F��g>��~.�4Ӫo��	G��XC�'b#��,�+4�9��!L��kG���7��-��V�Nyf%�����K� �s�Wl�q]�{�2�Q��D�~�;���)�P�ܑzI��4�oK�/��Ġ|�֕׌l��q]�EgOhi�X�ƫ�V��_Hf�BZ�.ŗU�>����ǡ�u"*eY�]�L_RQc�J2@TP%d
s�rj��� D�����h���6����5q2�Fa�)�@�t��5����.��f�����;�q\Y��'���)��B#R��%����c2�QU�g�lklQ�����Eaq��V�$����e��,��6V`A.�?+%��<��}QX�@�ډv"��/��9D�8�U[�&��O�qN')a_�ڛ�,�~K%�$��LEN���Ltt檯�����O�:\��E
��o���]�62V~@X����k���pPk�ֺ� $�5aJ�7_��q��8�.
���@�U�����)�iZ��6՘=��ۚ��{�?��A����ׁ���gVՑ����!���=J+�����k{�D ib�:TGe�����-L�[?�N����	�8��A������T��7�>��.v���>sGu�"Z�Ҏs �W鯤��!���uf׹R��b��ЇS������^�^U*Ʀ����f�c:.|������Bz�[�C��Z__VE�H�Cb�=h�b���D��M̻�JJ�l�*玕XN]�D�JŦq�3-�Ҩ&<?�0��v��s���xĖ�/�0��čz�#��W��R�^�'�vlm>|eB��0���@*KTԧ�Q �!�Ĩ?ୈ$}����}����a����0T5A�v���)w�{�8)�͂�#S:�~$;f_7n��U��]�0E�t�Ҋ���F���)U���>�WGY��N�k�yk��#���:�0���o81 �5�,%�p�E�F��I����^���Ώ���co��>\{=B7�8���B��vg�wO���	��1*���=�-Zw	����>�n��sG���|�x���,�đP�;��S�A�i~zUI����>m&n�H]Ru�"��[�;R@頫E�)-F�V,�?�	��w����őȚ\�ቯ�{t�f���h�4����/�X�r���Z��Dp�4�Qė��}�r��çq܁^
]w�f�h�8u�{���#�d7*ϲƦ&�h�/ l���k�/�Q~����|�(�P�I-��� jB4e�굛|>V`G:��
�6d���H��r�d����9�$(؉����2�3B��xn�Ѐތ���f�������ξnʚm����i4tUYg�~J6��դ��.�?����n��Sr��$!��f��8:!^�{7y$â�=��*������-VL<a#�i�Fw1c]E���B{��|�3�X���"Bz>���{�L}�h�f�&���L4~'q+#�m�1�e��{���� !<��O]�TJVx�b��bXlxVHYEB    8c0a    1480[/��J���o\K��c�؃P5�aᰓ#U���*�b�����xf�`�r�f�&E���}���K�U�)/�>ԅ�.`�she��!���{��	�I����2-��o����}-��.��}Ū�F/��a_�Gg%^�%����|!f
�a� �yA/��u0���p�1l�n�����-`П��z�O1��&����b9�;*1j�j���+���T��z�	��$G�b�.~D	���uu+h`�]��)� *t�iͬ{n�k��ĠO���*����ܕv&���ԦЁ�=�-�e�3`e�YbE�'s�R76��M-/;���[g>@r���դ�~�Љ���;�|A*l��Ёx׮"u��W����w��SB��_{׍TF�t֯�Iy"���W�ڽ=�L��~��A7k�3�䣤+Kۓ�����
Z(������ūm@��@�Y]zړ�L��L(�	W��aO4$�Ie�`ک5x+���U�/�{���
�5Z-��QHKGb=i��#�ܖ8��(�V����%	�+tF[�>�v������7��ab��e
��������s�)�m��IoE~v�{O�ެIsF�ֆ\0~��2b�R� ���c8���
���>]��kR��=ǣmU<�/��#y�T�S��'��!J�K�������l�O'8,zo>�78'��Et��U,��ٶa�	��$O�WH�Wcd9M\"��$S�Rd�����4�Lr�
���̝�������Ϊ)T�U �����	g�+���X�ѝp�)���oĨc�6y3�B-��V�lT�0�SN T���,�b8���!�k�Ƚ^�6"v�&�rz��G �l�*��K�� [��y�E{�*�����J���d�ss�*mF�s���R�mR�U��>�b�t���\o�դM��<��P/ю�������Ͼ�w�����&EƏ�n�n�J���
�b#�)�h��s���W);��z ��+53a�%� wo(|K��c�#�EU�s�JNfű�^�в� M�������4|F���&,�{.���Ƀ�+e�4��Ⱦ/���"�iΚ����s �ǯ�B�M/�	���|�}�d�p��w���_�>;�Mƚ�;��a�����4�7k���i2�E�߻\� @\R�~h��0
��tb��eg��������~f2������<)>�����8�~�Q�&D��^��E�o�@�ã�f*f3�(X1T�{4_���V�̜ؔ��bW��?p�`[�H�%�H�X�fˏW��H�	��-;y��P��a�]�_��96rx9AmV�Vb�a�S�^�������]/|�����!p��_U�	o8�	�¡ȠO���◌:<�y{������یB���x���+#E��/�P���K��/l�؛E���u!Q�۰@v:ްBM������M�%!R�
��X-��p�>f�&)�z��y�9��a�5�l�/��J�cP^=9�ѷ���豧Fm��&�x]�G��),�N�Z.�"�LJ�ZeQY[����?�T� �|����!����h��H��+4N~q���/��+g����Ulc��7�_b4��3��1�/�լ(	A���[��y`���h|���*0,S~�.���$# /�F`1�s���7�՜�p
�|\��ur�%���p��jj�Z�|)�sz�WhyE0�#�߾ф+Ħ���<Ҕ~K#� ���A��?�K'G�ޱW�@��d��0�4Q.�E�Ø�4���4������٘�L_��W*Pd �	)�t
2��ū!'S��}DC��m�ÄL,�̬�O!n[?��� B����ΡV@}�)�'�#F�S���٬C�����g	S�e�ue�q�������� 	�2тs�>&�F���XV�;�8^�G�C<�98ݻO&ס)w�q��$EY�2�����y���|����Κ!{�׈�~�C����ǮK��g3R	Kzs6���Y��r��rתR!'�����h�Ϫ��F4p� c�4 ,�W8���(-��O�,1�'����'�j�E⽩�.�X;D�A5D��u Ў`�����v�@z�hq���0�Vcw�3 �)�$������p��3:5���-��KUN��t�tn�&�33�;���[`�pw��n3C5|�E4�B�w��z :!���-�f�m����\�ܼ�p�����Mʩ�a��A�ޣ�n���
T`��b�'�k�;{����7�e���ۊA��
@�����[��ʹ��V4��/�/gX�Fj�]4Y�.�V�CZ���-%lL�]Cs��c������k�M�>��RKd">=)Ss��j31r��Y�ߨܙ%��Y�fl�# \��1c�������x-_6�K���� =6���g��,�Kx�?�6l���Қ��D��|�˕��_P�V6�ҩ'�&�O�Ҹ����n�7�o핢���3���Z��;4<A�׬*�(�Q
�\u=����=�y���!Ƙq��y��	�7az8������0�Ǩn�&{Ǩ��*��H�C�r�X�t(M���7����$��ә��s~��n@����kfǵ�1����t��AM���ϼтn9m/S(gv#��yR��o�kb���iJ�X�P��
a���r7����(R�D�9�k�b�.�o'{�������-4�!/�ʛ���_���$##���{�a�$�:H��؋���!�,�����t���Rg���0��c�FI�LeC��7܆D�ab�'0��<7��I�X̑)��G#N�E39��f��`��	 �J`4X=kx/	n\�xz!��P����ʻ�c��,��M�+v:�,�zV,�7bV�"��@qf�1O�"�ϡ��C0�=ѣ�p��J��>
���X�:�v�%u`�&�ʱs� t5�q/`��[^�$�R���������%�H���N�k�	��&6���[�?9�\�F��H�Pe�1)���9q�e���>�͙5	:BS�SgL��۾��}?�6�^O������R�ch��y���p� D?_�k�i��袠��O�10V�\!	r��5�3�"W7bI����M{� ���T���&�3'���$U�!i����/����`�c���(�OP��������
������nE�p�JEE������T�sεNF�gX�J4�ނ)�����9�?��=�]S�Љ��U�����U��V����#d� �<hC�$����C��gȩ�7���[��m6+��r��R@�s����14��mKR�=�x������M��8�����vT�J���3ǘ�^�e*O�j�6{�0�%���զAq#c�m��(�*�Cm�8����ˮ�#Q���ۘ��:�f�p�3����s��4{�^'����aʜ��o`��0��kO��(� E��wP^�������I�.�9�ᐎ2���:�f�CQ�a~�'�i����dI�1_��_�U_w8�]7�����2[&�c���^���QR���}��!d�O� =t�v2O1�.�O��D�s���i��l�fn?�7N������$��h"�g�5�IC�j�+��ίD@;ٳYV���������/�ｯ}�%u�b��뛩�*ŋu�
��&ew�ā+F�Lu��*IT��?8����(s��8���Bh���N~���Q�
��V.8�MEdՏ��?�&�g���	��W����G0�z�Н�#�@=��/Y]����O[�m��>�ֹ��F[�M%ٓ
���h���BI�xj�]R�[�=<���1�2>H�$eN�H���ݚ]>-��-��0P{��'˹�D����BlF�/�T֐U�6�	�G�(j7�1l�u7��������¨ Z��|�F��s�l���R�x���/z� ��F%gY�Skvŷ~��,�[,wX�s��M���;{ʯ|܂_h����@r(�˱���h-��308#b��;�D���L@��O6��><��b����j���W<:f�O��� !�H�[�u��u��j�B��ON��m��o�
�)}���/��_e���"D�ُ��U��y3�Pݪ���Z/��`��!��C�*��̫�,�z�K4$�-�rK�)��T�:��j�r����"%����y�h��ط2R��y���g�P���(��rpc��jw��昀F���������Wl�f�f�L�z�n]�U�m� ��S�ٿm���n-ͨ�}Y��u<X��䳇iB�����14�>�0��w�{R��������yF�p־�iUl����f�����}��e±�kP�Ph/��pmdޚ1�s��y�.O���R}��%6Jc��2�Q_���6T�'^ݵ)`sê��('ܙ�ɲ%*�Ȕv�0'B� _FL�h2�F��*5ZJx��;�H ���`q0f|p��2��j4��QoK�*��3-d6�)S�xJ��m�:��FOv��X�PV���(����pw�A���98ǚ&�YE�}���Q:�St��_v�6'3����G��Y�
��8d��	ǃ�|��!C�7p�ytǿ��ML>2;<k̌t{�1�(y�����Ϝ������,X�~�/������c����;��$��:��˶��<�����G�M�	Z ���!HM�!	����=:�	�+���R�R
�
��{�2�}�>�غϯ<�Mn8��b�ރ�1<.�W�GXri�pg����5-��!�ы&{y���P|6�a�	4jUMgǒ �Z@ �Ta~�Yky�>�1Wg���T��/�=�P!�)��j���S�16v�"+ݞ�W� �2#��9cg��F����Vc77�n�ɣ�0��|Q�b7����[��˟�}w���w��;'n�z�g?�}5�~��	��3FT�.��C����V���` ��J;VU��('�Wo���W�¦��[���6;}�̩��9����X SC�j���C!�aд���$�ܗf2Z�Q(?�m�Je>����PN�{[�9����@Ei���V��c ����[�ˊ�L�p#��+c~��Ɇmf�	�������#�_6u�Jt��Hog�¹�d��$�/d
�� ��Fi�֔�%�o�U]{�D �П