XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����i�MȥKi�DԮ�UH��YA�:%a&cw��-T�Zl�L]_O�����+1��Rh	I(<���b(@\���(ʃ��)�#\V��e�|G�ϨV�F&��J�Xzaʡqj�7.BUq5�d��;��\ �;uG���P׬A�L��/�БI��!_����ǃE�cd���%�`n��vN9���|���|WM��ֶ$�h��l伙bӼh�~t�q���M��dx�w��&\a�_�e�?�aU�X.R�\�YPʡ�>G�������ݧ�d2b̮�ɒ0J�Fwf�q��Ge�	F���ح��Qb��r��@�&}�`�E��������̼��� �,yFH�#��jN��R��8��J�x4iڶ��� �[�Ӏ�f��ę���wP����<���'}'?���w���"����V���A��F���	�R+��Pk�P���,7�M�.���0Y��;�	q��c�u�=Yyx�P�)��[�WC�v�{c��W�_·S~ł���.�8���$,sS����j���YP���x�ػ��\���A����9My�W��X�����ʨ�؟�m������#m�s�<����Ί��[:���{
7!$�\8�����Տ��U�0�	��iˑR�6�v@�}3M1n5� ��}qX��;Ղ}��ZGc�ؗ�[�E��%^������C?˨�؛ ��P�
*\5��T��kc��]T�����X����Iɮ�y5��	=�"ZWs���L���FXlxVHYEB    9a4c    2f70K�<}��{I3o�����{�i�-Q�-���.��z++��܀.!86]#[Ⱦ�7��S)T�i�6�_��jk�9�X�Id���Q!����)	'Iykf���s����;�ڏز�%q�)GR	c.F�O����X�(��W����7����ԯ&�+�7�	Agy�>����0B��C���AM�J��;�>ufKV3�j,D5��1��6@���l��6��ғC@�)~uP���GU�p^��DT�`.���:���Y]��"M���Y��g���Rf%W�hK̨%�ݚ�#�K"��:�Q�vf?�E����#�`3Mu����N��!�+h�,��q5p�~�)N��K]O�_:c'3��+RR9Ӱ���t[�ݔ�ޝ�86�r�~Jk�E����)�(��p�3��2+:�L�y��ѯ��̡�ƍ`skϧE���ѤӐ�p���
���5�Z�פ_sY%�0�H��(fm��p����;a��w�X)���]���?jv=�(�<y����M0��rB|s2%�͆��%4)�Q}eQhqC��w�"|�oL�ÌV2��e��C[�!�q�B#&��O&���=s���o��a<n�Jq�]��r���"Pdy4��΃�[-��:~��`]?�E���a����&���~��o��z)WdJ@��M�N��F��V)g��B�쟣)�O��	�+?�E�|���1�[}^��p�>sٓKY�g�[�G�F�lѯ֨[��G�`(Jg͍�VK�����;���(z׸T��H����¤!��Zb�.@�+P���R^��xKDMU�Zڎ�����J5�J7����:$���&γ��'����Qw�扞J	'j��JdҴ��#>���\%�N�O@x7��p�?v�#THD�*dc\���;>��Wz�<cg|ڄ�ӌ�Ƃ���a�$���� `��|n���W�U��t�d(7�TƔ؀INۤ<��sc�ts�X��J8��&���^�X��Vn�TZ(��d��uA�<�Ȕ�18�7�e�!J>b��}���-H�Se�e�7�M�Q������4y�蹨�.&|a_O-`����|�8:v�\��17Vf3���Gb]:�<j��o-��I��@�ueL�?wU�������@������9�E�e��x=�l6ÁƢ����y�A�Gy�l����*U����f��H<�!�E�߾eQ�Y�c���Ku�~ `E�)�emC�M(B����gDl:)T��)r#�X��e�2��6LTx�1w������:�>mas"\�C取�1��@�~��	�6Pl�t�sqx�(��X�^��8��.���i3`
�G��:�q�A%���[.�xq.����6m�f�Ydb���?P�X�_�>�k�h�<}MS=�����T�~�yWT��=����?�Ѓn��E�f)F��:ղ/�ӊ�b��k�7��xa�<O}n����*�4��U9�8���گ��Rw��L�T  l!�]SA-�?��O/ڿ����t�BQ��ץ��Hb�x<�е�"U�"`������P0��sN���-
)fke���Ԍ`f3���>M��m�l�FY�и�DE�$Q��b�qڻ%��D�:"
(~��L�����t�g��+8~�V��6;������o�����l�䕧l�?3�E&�L�):\���Ж��[���!�/�)�|��ݸx� �7I��`5�}���pfՖ�?0@�,�`��9x��<6��Ɇ����MN�}�%�_q�V�-��������G\&y�N_o'����B����j��|d6�tY�ʳlc��r�$B�?�a�_�?��la�f:��+?o8�3uh�$��\K��!"?Tw�Y8V��Ĳ���g��8Q���*vҀ����nM�i��f�T8x�n�ōR%M��A�}��*i+���fP��IN�����p������~��d~�Nؒ0v��>_��V��e\U7��ն�����y�9�x lB5l�}ּ�1֖	�U��� ����/FD#h��V�D����rǗ0�(�x"��J��*Ƙ5
��m�'���l�/7�Ri6����;���M�{�B��Ȱ�߫@��0*�Sc��[�֩'r�Dd�a?jT6�c�c�b�4�0�:L|A�:؀[B��I��$� �,)@И{����#$" �U��Y4п ��PD��(�Eo�c��D7�o����+�i�z[�>�̎`t�¬M���v�6���Bh��%�V;� \2��  _�qm�K��©�/�=�L��0s8,>�r�1��HF�G�O��EA�Y*ڤ��㉎��oz��e讋���V���E+,��$�d��ϣ�:W��`(���S;́&�[��y8gO�JύF`x���&y��n(��L�����?b�RF[�����F8w��+���Q7��=�+���'����`���`�����_�Ѫ�P�)�Gx����?;D�hA�"�+l�L
�kY�*�N�m���^����L���@�S\j'���
�����PD������8�f*卾��H�2�Ƽ�˨K��A��y�`���L|���K��&�e*��X�b��7%_��1��E�D��b��� f�7�i�|�U𒩃�N��:��0�Ep���S!�:#u��ޠ�
�D��I
�>Ldߚ�m0GzSI���L|yC��_g.���H񊗳�)��6�C�}:�//G�ꯂ��Z���?6'������gf��RS��N�]�uw.a�Ze���c$���|6��׆�J��'u� �I��ަX�)���eD	|LDU��͑���p����$'�[V��|����2oNr^*2!�Ѫ9�Aj��kV"��M��[����&�̀R��V'6��Ih��F��V;u��Cǧ�U��2,�q�"Ѿ<D�` ����/��J祷lKG8J�Yz�V��ƫ��[���6Cr�����y�8t����.����a:S��7������ǧ�	�t��L,Z��:[�9��;�R�#ϺI�4�l0)�vvt~���2	)��E1c�����L��}���a��/+dR��kos����#��`v�����6D�l�B��+9�6z4�P�;��85~��e���{鍭	�
꣚̈́:�a���/�*Lx�7l��=�ϗ7JD�B�d���Q�xEi��\�왾�ոڕ=i��w�T�|�2X�蚍D��4g�ȿ��ݻ���Ě���[\��@�ͻ1N�=x��W��_q�였��%V8�����>��Cf�����>�"0�a@ �
��p�F�9�+sPG����$w�?��bz"�8����z.V�M��T��04���!~1q�u\O��/�͒��ݫx[�|dKi��a�>��$�����n~�5^0�1��HI�&݇(Y�r����1��s�d��(�A��(a�_^l�����ě�5���"�oC�}8e1n���$p(�x<gUW^��U�ed�۶KHF�� �qzGF���˕���mפC���>���6������a��;�*����ሚL��R�	3VyN��%ѷv-F �'v�)' eQ������䆊�>T���˺W���_���U�g{Ke�ܐ�<�F���V��FH.C���~�wJ�,O֎��c}w�%�Pѽ��ǰ<�)쐁�}-A�,6�JŃ��^P�� �{t�
�/q\��f��k^��W��h",�o��� Tc���Z(�����L�7�	�r~Ċb�:n�N����&���N,N������OH	܉����06��~�$Z,�"ѭ�V����:�
�%���T��W��u����3/����c�&�L��Aj��P� ��أ�My�V���ɟ�^[D��=n���2�ɸ;P+�>^���Sj{�f�d�V�4�L h�.�2&�A�0V�g�Wy����x��uf���/�]p�wg�K*W��~��B�V���c{�N��Y;T�B��s�>FY��*[j����v�*�E2�'��Ї[#��q�6�X�SJ�����^dٶ�s8�|Pe�N����Nz��J�)A3�G�@0�Sy6/�e�m�Q��¼j�W�a������9��@��j��� �(���T�Ab @kq���,�2w�5.~1@w#�V��T,ƣ?�����`�~%�;���偓���R��?��7���aL�Ce�ٚ��n�s$�R�a����#��X�ѪnL�^@?9���._l�2!`���0j���o��ApυJ_������̴���Ş���)&,���5s^�[EC�W�J:�yt$��-�}��"�Gb�g{��F{+\t�[X5I����-i�0{�w�:����,������^l&�ܳr���]H?�\�%�r���HΐεL.O<�W~���� ����IVo����D�p��l,���vQ���҈�[1^�F�]lI%Lvp.-,"��D&r�f~4M�b����m��	;x���҃������B;�D�
�����
�����&�X�c8~�������4zV�'�{����a\�-ډ�ܺVɎ����|6��k]�5��$*�����NS
���/�{�Eo�[��A�
)	����I����7PnЍ�E��W¡����F�6��?)�Gq<I 5�إ�@T`a���+
lf[��#��m��쮻����l��:6����ǌ� 8[BmA�t 9��T�`	Y���y�w�*ԎO����MB�x��.:h�a�Jx"HgC$INp�nҗ����0�z}<K�y�]����H��5�d�2a}{����v���}�� $�H�:�ZǁX=u8���f�3�����h.ܰ�6��^���z"}Fr��N)��6���?�8�3HXԣa�u�.3�d���[Vd�t��f:��-�HB�0A��ݤ��R�WO!�ؚ�{�+��@)+�|�e�hP�S(��6���J³�b�$��n����*�G���t�%��EB�9pN��r���]|ݫ�.�Lb;�E&���IK۳���"�����Y}QX�����hL�_z��N��"{�:9��8�Yܖd,�zm�����;��D��KW2v��?�PGY���W�!S�s��w-~��p-�8H���qa�X�-~p{��|_�i�ص*��ܚ�"��Gb�b�����̨>��v e�wq��􁑍$���)�/�e*�ϣ���u�y	����/�3�~��L^0Ro�}�͈)�
���569�	\��	�Tx��OA)"���,tWg��	$-I���*!?���w�б?�8@��ǹ^�ڼxI�6�OQw��޹�ŭ�,z��ø%����$����lt��wI$8a���C:�Z=ߊ6�*������ے�5��n{٦�G�W.CJ�����q���(��2�����s�[R 
�����4�$Ē �f���0F��C��Y��=9ۦg;�������֝rt:Dcg�>U�P&:��:i \���m^�q�U���`���$ʙ�?>�Z��V�L{�S��E� ���߯�J��j׫�/�ر��J�Ǳ�ii��+ߧ�f8֝� �M�3�	8�`Fa(��?��ȯW7���(�X�h爙�b�L��@�s�ˋ)�@�N�n�	�aJ�j���� "a=�`�nr�e���R.�_��	KVv���ŬHh?��h���hr.�t��[����������]<�)!�2y�������K�І]1Zlom�;�=�Š��p��AaN=�v�A��2	�{�1K��/��%ӊ�&x�b{e�`\�qc�"`�A�_��:C^�gԞ���wz�Z�)����i���K���"����S(W
����@�u�3�P�/�����#	��uo�|��w�P�A�T��y�b[˟�:�`���ΝW��!��e�N�S@���w�\�׬�2�3�d���d�^Ge�GMd�F���N�10ʠ���FE9C���E�Wϰ�GVG����"��1�ϟc��>�:l�B�//X$�9����TB�
K�����<����'%��<�J��k�A�j�VR�BZ[�[���?�&�㦨��L�-w9gV�� [��L`�+�c�;��!4B)�������W:B�m�@�
�t#�[<o����֘�VoC+A���Q����p�@?�9���vTZ9
j�W� {���C����O���*-U&���K$.�=_���G����_°H��q`�� v7cU�Wx� ���=���T����f�H;�$�g�Uj����D|!�*��i���4�?l繫r�`����Wչ�(�fZ��n�k{IO�� ����6ZS`YY�~2��K�e1�k�0*D��<o"����k��@�uC�W��B�.���a���*Fl�C,�Z�ԝ�ʽk]G�Z�P��
�I��r�A�F�^�)�C���R��@��ϱ&��ZP���W�������srD��5p*��ۅ������Ŧ��1%���0��hߠ՜9�(�k�;�C�z�Ŭ�q��g���I�\+D$�[i�N4�梙�#5�`Ǚ����d��4�$����k��&�F�(Vd��@�&����������I�;��L"h�k�Zo�j�3����!�������ʛ�8���Vv�ā�#����=#jA^���#x�i,�^8��UQB����h���S����@%v����e�j���D��7��W;�eHy}�z��ohj\
OX��w��\a�7�&�H�6	9_�J!�l��~��S���3�=��9��|��P0wa3��A��$z��t�^g*R3n4X��]Y��e4u�e�c�.w�m%T���n�Fӽ�W&Q+����UH��m�,o?�
�Y�z�*������Pe$oМ�O��;�]�lR�FW�u�M[�}r�(/��FS7S��d�fq��\���"qu/��ޝ<X<�q�#a6JX�2�[�'A��+�{k)b�,'��n���EY�m�23<�ю<j�h_z�q� /����z��K3 x�&��\|!)e�����-B,��`%	�0߻y��W����SgRz �̿������ �tO��w�����u���o�+o�4�/������ҿ=r����Q{>Όx�~S[��ũl�`�*}�f�|�W��P)�J5do��t�e;�Ķ����_q�%�\��w9��V�~��]jX�O���V��q�LԢ��q��j޾��tuڰ��������'p�a��xð幹��kOb�c�Uq6������q�	1ڄU��x5)�f�U��ޚ;H������������X@�� }(�.A)�AbԢw4	ׯ���/	�8�c�ܢ==�rQ���/�QS ����s�����*�Ej���g���u��h�]�~_�2}������UU���~;z��SA69�N@��K8:qb	�2���WM&��9c��?w�h��[�H���y�¥9�m�c��j7�}����5Xc��7�'*���U����N��v�e疫I2޺��n��j��t`�"	8՗���>�����0ż�;�eY7�������'���8��N �5dFt�g~�#Tqm0p�
���ZJo\��gA������.��k�g
Q]�?.�{�u�S�cܚ`����޲jW�Uk��G{2��c�q��֫R;���/]�"!9������c�^��_ʍ�z���/G�wm5��x�+2�	-���f��x$5�\�#�}��8��d'��C�7�H<m��	�CӪ���w8�I��@�|n���:���iͷ�q�zՊ�!!�9y�5����6r�� ��׬zԺ6"&(Cg��H��j��D��g�ֳ𔦃5~���>�d�
���5��y�ZElŶpD��]�<pOu��{��{�*��3�eވ���Oi%{7(�٫���qz�ʜߜǏ���0Tʇ�'��,�=��4Z<�@?8�T�qL0��+:���<x8_�b��)��;Ɯa5�P�ߟ���X�>v=ާ �ռP)M}� n`���H�1�������R��g�qJ��|��P�>h��"�9�4X(G׿�����_҂u���h���])�)
�4��[~ؓk�%"����2{j]�̘�Z�	W��R)Q�b\1 A�
���%L�z�1�3�H�~L���ޒ�Ynv�Q�z�D�x9��Z��,G�q�U��b*�7�#=���o�ĩ#�~�){"^}-G����P���Y�l<9�y��}ti'�8:I�[P䉩DIp�8�O���ݕh&�Bz�P��=��ɟc��>��*ТyFo����;U�\��NS�u]h��|G?�+�_y���&��y ��X�Z1Kn��Ny��	upñB�ϑ��w�3Q�Cyc��-}�
��\��|u�e�L#�����,�ս3EO��]\�թR5���T8(q����v��yd�E��V�I��-�R�8�AD,sb�B>݁L��g_���}Tt
n����b��N��b%lm��z�R�SLJ"�=q��K������d���Τ�)gz��98�c0r�'B%餤��|�L���ᒀXd
?���Bߪ�,��P�����m өE_+$ǐC]oG��Ųi�^�Š�ۗ�����nb��Ӈ��b�u1����CE��� ���j� ��g�:�2��PTk�%Ek�8�ր�$�vϯ��l^��b��^�!~���ֶ	��N�K�-_`��!���Y f�! 5�i�Rq��}ѳP��X���V�����;����}U�c7��CU-���NG�F�"
����Jz���CC�$��v�D	�:�YvD~iՈ�C�r�=쏌��s.ڲ���P�9"���� ������p$�����C�yK �DS�̈a'_�}E�������&��ˬ9�Cr�EL�:���k}]�R`}��n��0���Y�Y�Ƚ�2.oX���w�QN�3`�$<����ߕ������k;�2�C�]��o^�(%�V�qĮ� �ڰ^�s;v���Gl��MvE�@�e7>���/����)xP�h���:^h�C��V*N�LF�L��^,�V��hM�6��9�Ek�"B!bX��HB+`
��k��������ƺ��� �����z��[��:!yڄ����K��Ox�*[��zC>��F8oE��JL��hԸ$칌�l^goZ��US�\ۨǳ}��+*���k�q���DjM���Ѷ<j��D�m�+��'���2%(�����qsD7�F^k�p�w��*��_|D�&VR\�1DS1�U'�4/��tS�����T���d�G�N-�������J�r+����Q��nkZH�)�ʼ�� wF�\�w	`&��i��8��Glm?��@���ӟ<ˀ*?Z��?	[��#\����lm���T�'��R۬$E�h �E����>h�d{Fi�b�L�n���1������	i޷2�[��߿���f�0{4�(H��I��+�n�}����o�1�����\P�y?,*X����wXy͛��ˇ�SwoYLz��]��\!��[t���D�?5;8EG 	��2�_�D��r���>s�\u0�Xݝ�^x��K3�E�C��'MM�QE���<�yRȰRg�{�[��(b[#"�K��B�|jGr֣;f)`��Y������|��6�{�� A��<}�e�'��{���Zҕs�0��ÆRR�4�Ic�a��&j�j8�]T�K\�術���l9Y��S���g��g��x�>�4Q�"����e��.�4��\��q'\���g/ӽ���`v���/t�<M\��Z<cSY)�P�uR�7�&p;jC��s��+���Ic�@�;u�q�|%�BJe\:��ԁ��\�A�}n��Ͷ��y�R��aM�`��(�v��jkA�sG�b���R��Q��m}���#�˖~(M.��h	k[ʳws"����Z�v$&с�_�|'�!�qLC[9c?�xp^��6oi��^/�^����bv�ܥ+�x&��AD�������4.>�u	#�rU������Oie���J кv���Q��z��g���dmet�Ƭ�&��9��4��ŧ������7 S_�o8�zR�S-�(�a/hٙWo�M�%��,7k�s5�E���V�1��=����؛9��9g(�X7c�B���<~|"�l����Z� �99圍�+D�zA!EW-��G���]����g�)M�Y?����r��,r�v��ҋ����*���M��ҡT��b���Q��-��_x�I�͞�l�|r:}�d"0�*�����G3G|��Ҕ��oH�~� 6�($/X��a5�Ǉ
p((�]��s�D���U^��ُ�Y�����dM���Kyo��y�c5�G�v��K�F��/4�y˔�	�i�+J~�q������I!χ1�鸻� ��H�8�r���d?EX<��ֿ�6�L'���A����y-GI ���WN�z3�� �����{��|���1s����	ݮ3/�Yb�2��;��tOQ" ����O2�������瑆Đc
�yzҋ��v�j�4[	�O��q��6LL߅�^<�U�>Q���Y���v�a��SNlE"jͣ�fD���4\�����]
{Ў� k��"��?�ޔ?�@AL�:�"k[ �"���XEǂ���y��R�JsvUׁ5� kp���cP��CR�8/�0E#�/)��Bl�N�lzAl�4M��\S��G`�%At�xyփ0�O.X���"�}|�'�%�Є���|�Cі�%�܁�i���*ʫ�u7v�	�C+i����)U���V���=.�� ^�)�9��8ڦW"�Y ���<�g�(@&)LM��'��c9�l��{'���&��;��RJKA�$҆nD� qn�A岰��q���eX��v��*`���
�x��VD�=�h��_�P�
SD� �����>N[)�NN����k67HZ��p�*a7�	Q>�)�m�Dv���B� /K�f�u5�a�[ˬ�C��<-���8K�3��Q������{=j����f}|�6�T)��C�YM�R��`���M>�gq#~�=Ax.�hCҗ�p�wFq���h�M��$Ւ��v���3��1#6Ԧ�4Kf�ͽr�&##I*n���z�����u>�2!�묧�\������6�Ҝ�.�C�/���`�cK�-Q�]��ō��TM�ÜN�MK�HP���[��%�!���}C�#zj��z�ܤ!��{X�1@4�~B�+F�o�M�t
y�%�� ů"&jJ/t�����v��K�kGKO? X�is�_8�C_��ȥý��_�o�/1�+� d1��.r7�*+��8�9�Gј��;�,�Ju�V�D��}$��cY`G���tޛB��r.��ȏ���V�'������j���t�{C�si�b&�io��jQx$��HJ,��c4*:'��C��=�U���Z�o)�C����3;c����yBbE%	)C <�%/8٣�H�'�����*����f˷a�ʏK�V�y�#������|r��b�"f*�A"ƚ�Z.A�}+ƞ�<f���	^��vn�[^�d���E�H#������&�5~
[��.�Z�c�ʵDCM+�ڟ��kN���#��('���_BhE��v8�D�RB`��͉[�B��XT+�?�p����p	ϰN@��>3�m.�5f���髐��u������psWȖSٍ�5#��$)L�C���c�-m><�z<�j�����[�Y�%k��m�aZ`lQ���˻�vW�ka܃�2�&<'Ȫ�Di�4�8��3����&�e�Y�i[���������Թ�Q%(|0����b���	������.�/6���
`�~�>�����#�a��	�*<ɷ��N�n�+�