XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C����L�Fe�,ʗ�b��(�HN�8rgٴ������ţ�,b΋��@�%��`�
��s����@C�)��6��xئG�>�6��:ep�V��@b��T5H����(A����Zo6\��HD��B���S�j����
������
�S7Ś��ZF�z��:{h�/I��ܣ�D:�W*��I���GQ�1Q�[��D�ע��!Sᝌ���v�A�p$+H��8r��+�����r�R=U��h���3k����1R�2�l��g����<��G!<2Y��qG^�t�ꂿ_y�!����׶6�1~�ͬt`����6;�V��,�۬6�Cu��P�a���Y�����f�^��:�!�������{�
���5���&���t�7H
�9��0əX�^q,�}�^_j ��UKq��3�4A}���`�
h��x�?0�~f5��Dl��j����<E�=�P ��h�����ư��"�P����-��B�b��+���ֆ���Bfg��!���+���E���ݞ�[?�z(gx��l휡K� ؖn>�X<u����qO�_�I�pY����W�9uq����Y?�뿤���|%�BA�Xx�	����2"C����aC#]�ɑ���yGm�� 
�ӵ;��r�x��e��@C���;;z��)�Si���_v1�'��{��¶�E�$����y�\�Z̸lx�Kzr�Df�HD�G[:���u)H�~��zф~l�iw��XlxVHYEB    fa00    2010���t6��&�h��q,��j�w�j����D�K�J��"(u4rn5�b�Ig�8�b�Od�Į�IVx�t�xQE��!a��7\i^ョ�p��r�)�༯� ���Z�xḱn���VY���s6��蛭�0}\��9Z�14Re/�;<0��f�C2��r��"!A;ж�����bm����|3�tJJ���um��Ep���ܲ�\v��h���S�hi� :�t��U|��[�Œd�4
�&Ek�d�p�^z�H��^�}VJ���\�+h�
i_��X�G�ٳ�/!*7�ynZ�dI�b�4T�c��@�y$�x�_��B\����	57˺ֶ�?���:fE�S�W@�(;��܄���Š"�����[z�-����)���S" Vn;�h>���h�ƀS\���&�)�=�Ӷ2N�%�ȩfâ��oA����b��žQ�)�'�Ry�}��L�yĬv	^!uT�f/Goy��^�Y�i��,�����!�����AWeR��H��M'�t�����f�v��������Ɗo�4��G^�|Lq��-��K���3���Q2M���9��W�ـ��P�ؾ}��bC�|u��8$p0�'��n`��+fu��޽!��0���-T�8d���0&/�y�v��U�K�i$��ӛ�;�ԗ�2��"#0˔�8��v��^�TX����.= �Jj.�T�UE��`���,|{LQ�a1jU��1Y�G�u���Ur�9{����+|��f�H��n|t���}������\/�z!���9�VH�T�q,��v.����l�iKZCu�:���)]���]����b���X~�,�B=������=I�����Qp{u����0�2m$���N��LΖ)�ua1�C�o�I������r>,���W���V�h��4�o��.I��Ii�`G��N�TyK/v��v�8�ϱ���Z2\:7������?�@�iK��#�J+�		�h�d<����B��s��ԑ��0����5\�L����N��#?���:�Q�̶�ש<��c��G����#��*��vu��,f��1�nO�Wֹ�-ܩĈ��E��2�~��#��#�21���J�wR�Sx8͵~D�sއ�/K�0C�Q[wO(t�ť�`�D5	�}�g:�Qk��zQs���y��{nr�����-ML�a��&o�ᓱ�$����Q���67���bsԱ�����e~Ԅ���o������y�]�T�j2w�T3��o�J�-�V�r��/����w��� 4ѷ���1g�I�����bT����0qQ�%�z�k�����*�� Է"�&NU{h�:IY�ɴ���_�-��&�L빸�����F���ox�h�� $ިΧ}zD���z��{p���B�4�K��P^(���'|6p�辡��� �=ה3��/�65�a���y���勩Ԭ�F��uV�/�+�
�-�9Fǥ�4]7�w�.6�TR��f�6�$���Q�<PC�FDug[��>�!6��Y�
��<�j���E�t���ٿ��]�mp��O_N+s�8��PK&����ŷ��.���|��常���X�#��Z�s`��}Ng���.�{<'����h1��dt����ZHc����[kRO���N���B����@	}�B��!e4	�Q�L���cm�W���c:���d�� nN��nW�u��
�K��΂�!����=Y�-�ߩ�/iY��I�����g����	�ׁ��d�V�C?Pn{�MZ�gcQ�.�V�}��Ņ)f�������,�x�V2va�W#3�jI#d�>aD�2l�b�������ex��'5�	-���0]���b�V���{���;BQ���� Ð�D�Ǩ38��&,�C׎���wz{@��?�"%ζ�z%k��^��e�O�K�� *ҡ}'�L��P�&,b�Ĉ�@onV 0������m���8�p��q�����&��Z�����b$�k�F|�ɉ��M�����	d�ғ�=����0<��4M�wА[0��� ��ԃ�ո����o�/�������A[G�4�	���)H�OB��2L�,�]�`&����R0��-M7T�D�r�Ye��ȹd9v����2ej�#A��׍ݙ�K%��� �j+�^+�'_�*Ӟ$z5>�Y���~���!\ʥ�TZ�P�=�"`A\�r��Q�s���:�,�����%�<ZfN9�Q��n��Uj��_O_�1�I�"y!���:��i:��ӻ4�08�[��*�j�BN�ň���s4]<~/��CGՃ��nz��;��V�!�l�"��G�g�N����t`���lnLb;K!��W��hxe.0�Qs�o$�d��$�Q��5��~��f��	�{���`6���p:�|�PD�}�xh������A+>'��M6��5�$uO�6�T��-(�,�����oR�U����|����7Μ8�~K��N��(����$���3�]�7��5kZ���IA�X4{Se"x����/I�5��
��Ngx,4��`����.G]����
�Bo��%_��o�\�\1�Q�c�`���7u!]�6�H��Ic���7
3��wܑ�h9�L{���~��ܗ�iߝɳŧ������ގ�9Dz-5�/��
�����U�U��K��$�O��L��h���.	�փ�(#���Jd>��vy�q�5�mZ��Z�4m�7d���i*����Jt"Z�Tl����l�8�����!�Y��r����~IL��',�[l��,����R�%�����i�A��,˿��#@	��&9�9�iK�������V�ţ�|�q���'��x)�5xo�x	��@��i!)����~��GE�ak=��J��ĂӮ��u/qb�
�O��ᗗ�c�Ŏ�}2�狈�ڏU���<?��Ś+��Y���c�`D'>�K���$�*�;Md�&y4�U];$��F�X��Zx���"�o�늿�Մ��$�`�5M��$�"g�벼�"�@�	g���xCoCF�%�ӾG�z��h��xi�Χ�7if��R��&��M������/�)s����?���$�9AK� �X?T��$��k�Uj�w9gn�8��c�!Fl��J%>�pH�/��K@�����``�	��t�1ʣ���o���2U�<{@lkc�YB�N�������Z�LV����w"3�E,n4+������ZU��D�6QMJ��%�E.<��J��s�>�a.���<�v��Hnؗ�O�?l�;j�\̯�Ӻy/bj#Ԁ���[��<�(�� �+#;�E;�o�)cߛ5���؈��8T�����Y�V���
Y�U�g7��T���e��q�bl�g��������g�>_�qӡAM��0x$�b=+�n��ÿ�����p뻚�e�A6���.=��7k�'��@3��H�^���y3��v~~N:=��N=pd���fz��X (<�>"���g^����aݺ��VӞ���YA1Q�x�3��F�Ǆ�p� º�̠?~�i�(�e�Ks~�w��h���p��Ԣ�D�f�J?�N�"<V���tb:��#�R�K5t�%r�L\�s���дX9�0�ߗ��+HB� f�(>��*q�o�q���1;hk��x{��P3C�I{�c�(;I�VK��}���ة'�E�rx�:�0M�L&���EF(y���y߳�wrjl�cYA��������z|e�36�`�+\��ev{�0I�b�#��wZϲw�)��N�C��/O0[}��pY1>a��,��l��Q��ZT�<�)�x�R\s���� 90�^��|��grd�Z�Oo���-��g>a���i���ت�� ���!1&{�>������Xq:/m�*	�D�82�����7D7J7����N���bΒ�h���O�m�μGz+ti>'��� w�kF�Peo"�v�.K�����ǝ�I]�y�C�aJd�EN�
j� t�zic��w�Va�4�5�6�(B���B�|2�yQ�M�3(�xkT�s|^~
E�C���>�]���`�Et�#�Ji�)�H�l�);ƅ��X3��J�� �(w4�Z]�,S�e����ٵ�;��o2�w1�։-���#"�^�����m���	��_�f�Jw���@��˹+#jt�B��ږX�%�	d�ڼRN�O7�Mt�>v����g�C����t���Z�t�H��5���1�lܓv:ۏ�G��f7E��V�`��Ba�l�GᓯW���	��b%0$6~NI��B��C���Z�u\��P-ޛ��2g R��j����Ư�Sc���ȉ��~q��:M�,��o'9=�=�R$���'��0��n�09n�����֧��9�.I/*�	6�=���������Ē� ����<ibMJ��+=�卪i��ꥶA�kɓ�XhtNZ�2L�Qf�g`T/��i�<l���C@�F����-/�/I{cm�3%��{�|Z��rt2؎z7�/�{Y���t �@������uw�5G�{��\ZxL�jfo_px<T{���lZ�ӿg�UXZY�L�����e�À�)ߤ��1�����������T�Z_�KKEjO$�린Q�D�1�$�C�|���$Ք�\�,�0H0L���Q}�	8��#�[�%�jᴄ��@���(v�
�4�}'��>��Hg	V]J2Y�3V��%��!L(�W��8��u��5�M�m[)R�X��}��s��n䱌5� ]K�9�:�^�n6�M�TD*z�N^G-os��b@�ױ�{0�3+��SU�}������LtCפZ��g�o����>��j1Dl�-���o��d^��T�� �F�e���Й��JT5��m༱|$���t� ��H�U���MU���H�g�����s�$���̈MG��YS���kr@1M\$-��bb���_�B-����4�����Э?J<@�C�p�%BXP\"����G����z��?K��͍�nl�Z����k(�}�\A���ڼ>�)�z�Ó��r��n̉��� $��~(ocsw	�&((v��Z[&er��f�c~�����1rj�f����I0B�IdN���z�p�H�~���w�6W��C=�o#��ȶEl�e��aO�Q@�Ũ�8�#ua���腔U/��CX����c����xr&N�a nb�S���"(�^>�i��t�ч�L�"����6r9��QŃTL�3���N��Q�'�8O�ZI��j&�k&�AD�������a�Ǵ�EU��ź���͙���n�;�eN.̺Ok��0���^l��KsN]�;�3��X��0R#;�#��C)>��sdN�M��[��"}[lU����r r�{�anݸ@� �hl�Ǟ>���n�/����)�a�YY�kl7S]/o<���6wz2ԓ�� EZ�����9��R�I:�ۚ����ի�Џ+�Ԝ�:Iw���!t�_T�JX�e�p�#�ׅ�2��|�,X�=�y��Sy�)~D92�}�/bҾ��+E��m�?f�S���m�e�� ����Qs���3P���Ao����8�"��p��(��Urs�������C�w�_:H�JOE��^�V*�9r5q���v��T
=NșH��N����m
��{K.��8��D��CM�&�O�{�iI�?2	�1����%��TF8v]��Qb$aw���L 뼾hzz�ŗ�4o|F|��7�&�A{��&$�}�@��o����y\�k<ƶtl-�!y���9Y�0#I#E�4�ɂ��Y,�Rv�D��@`EX�=h6�u�S>Ch�����[�~u0�����¹���25�>�3���W�S]ef[Ɇ�F���${1��c'��X�4z��BȮ����DMu��@��y5=*9t0�W�$��3<���p��;9h��۠�?`��X�QF3S;w)*����{	4h�����E��=9�k�
Lt�؁�p��	���5�/LN1s�����4�3BQ����,�J�OG]k�e�l��(����tS����`s+�8�����i����⒇�0����s�����|e˒Wm�#�	����_�e2�{�F���j3�}2�{C1o� �����tY�sb�ws�t�*�L�Z���S�	�8��粕��^JE��SI�ĝq@g�h���%�]�d��i)�~�0���!�c����m̱�д�Ў��Q�����Q��Q����Q�X1ƒtG��H�Q֨B�����(7�ʭ��(��S���(2ѵ9��'�n�o�m|Rf��� A�����-��Ԍ�SE���U���,�b��u�T����D����,��2@����6ʓEi1��OL��"*{,R7��e�XP]���[O���������Z܎�6%�;�<��b����Q��/~շ3>2��_vD���Wi �5�+�t��{�2~!>�=�}�3-xS�~��9��Ͽ�IB?
}��
���Ư}��Y��"xLp���=�rA���u�r.eߡ
b����t��U�]Gj���e�#���\���^Ĝ��4���c��.Sp����
�3ǥ�?�ް�b9�|�����FY��Q���+��'���t�Z��sm��|���-Yyc�c�,ǜV3`Hnƅ�+�)���^�X�I��Np�uBr���f�R)���w�x�w!���MS��[���CV�}Z�ڞ|C֝��js��p�0�w_��wi~�-�~��F���w}�"C�����Nާ����@r߂O������k�y9h?Q�^ݔ�'cOb����t��U��'U6ɞ{�P�D��f��9(s��a�6 8��UW�l�o�r�OG�ŉiu���۱IZ_�5�c�&jnsK� B֌	)��!6��H�X��΂���q��d���F���aR �E���:ͮ|<�_�t�x4)�>��);u�."���4�o=��������(x7��%���Ks v˲"$ۃ%��i��0���<��l:�����.z�$�w�(Hd�B������uc,�Dp�L�*�T���i�>����󱩅�wC���e��7ӥbB	�չ�U��~VZv"��B2G��ц�|;_�[{���Җ�㇢+7�J�1��^�di�h#ފ�'�>y��Yk=s��m:���=�80�^��n\��-�dLV"�`�/�$��Yo8Vo=�0����{�&_�mGзVy����cӱ�يOt�K�L���Р�H��Z"�_)��`.$F�$�h�9�����8��i6�T*ȣK��`m�sP��-�B�]�}��B��W�Ǝ��0c|q��l˨-�Śf��kG�p�a#((��	��/���Ѵ2����B�:ٵ��x}�ՌL�P,H�h;�$ d���){`Aw=�ؗ��,o+$�K9���;������K�����N�(z94����[֥�� �ɛ+6FW{[lK
mM;���1}.�d��;��,	~��.�gǘ7�fM�K�5��Oz�u�!�y���-�	hf��p��2�d2	��=M��v��ދ�r��3����Q���=��y���ϰ(���������Z�ey*1K�+Hs�&(�Dб&�������͆�Ai�3�o�r�z����,x�b/�]`ٶ��JH&x����Q�PG�Z�0�?W�@)��5�lǾ�<�b��D�����I>�����+�d4$cq���g,��^�δ9���,�#�|�_����GZ�ɶ:��X��z*Z�����u� �HzY�<isW���v��G�����j}F9�ȃPã0'�&j_\O�צ�ց��=~�4ZtK`Y�8z����9��M��P.�%��N�f!�6VRo��)�¾Y��v�D'V�tQ�R-�"��I D���o�&Q���c�0Y�n�B��{SV�P-�}�#i�m��^�c������;<L�#��ޕ�(�1v}�o��g{� CB1�TK|-f�K���r�a�P�;!&�?�r�w��|�.�
s0hzl4p}��<�=�<�ȏ�B�N��Α���c��,�!:�ǻ���
Ѕ/LO͢-x9K�T$ xXlxVHYEB    fa00     9106g�0(o��%)��Q�K8u�����_�`	:{y���J1l�29��?�h���ҟ/:�a�Ȏ1�7e:g/���ߐic�ùܶ�� �������<��FӋ�T��H'J�4�Ԅ��	�ul#��$�����|��}��(�(%b���ȵ�=g��,n��������6ު���G�r�N�#���-�r��i�N�Z�@?'�hm��~��d���2A�|P6o뚋ݺ
�G���vCRPF�{p�kjs1�m5Z���?�P��,�&%Lٶ�M3[[�Sƣj�P��&`���mrY��ٓ�:����Oo��9<��ob[)/�#ޠГ��K�M��4�o��fO"�2�z����U�!{�D��)�����~eS��v�<�w�����:y�M�ޟ�F-,���VT��
[�Mp�\Q;;s�B򵇤r��6��yJtY�s�ߒ�ĉ��~N��ڄjE�q?�����"�17�E��(b�/��9{f�,5{UMuN��5�+Wb����G-�a�����I'h1�v�T��` �����e�'�\����k�ϻ\�;3�m����d��RMߢC '�Z��� ����i�f�P���S�vAC�=a�=b�[��'I,�0�v��s��/��1#S��1
�l̘o ��rZ�Me���փq��8@�yYD��ncH��8��;�PH�IK�N_bU�] �>r.� ����[\��D��j�4�rjKG�sЁ����O_�:'�F��,�Ӄ{�O�1���~����u</�(�>��b{���N��C�x�x�����缋���&~��|����Pж�&LP�SS�;��Ώ��(���1!�5���t�3;��W�]�ݎ��Zx�*1�[����l��#H�\,b��_�e�hR$g{ZE�b��hD&77�J|����#����?�`��F�Iu����0Y����_Q
���9!P�L27?T"��e�1'�n�#�%��'�Í;�G��
�5����j�J?RJ0AT��vMx��,��U��h	
z_��wስ�Ղ�Y@������"�2���+5d�)�qS��6�пM^�4w(C��P���O�e ��Tx��C�޲�d7*�1��E4��J�Q_İ�Y������@�-p�i����|a�#������}#���!Ϡ�������e�ؔ�p�e(2���ZɃ�
��=��z��^�������!
�2ug ���t����KOV�Tu��L��ũ�O= �qm�|F	��;�~��j~Ʋ��c���-HC.'J���i�B� �Ӊ���W����d���p��o���)x�h^���2��C���˾@�C���R�&A��
��JnA
��e��2]��˅�r-XZ��F�f{�c8`�t����}lڏ�RjXU4�X�s�Z�W� ����i�"FR#����6hW��T�s���_ m|�P\�br9;%�]�����T^+��io[�ny6����UQ��Lq��P�5y�D�>�}��[�m����(4A�s�/x������|���͡YG*N}��׶&�O.Nx�7�h�&�y���wu�&ݢ̴Y��1���4ۘ~Y���卓EN��>J��Q��$�.�;�ݜ����]5�����qv��6B�m��UgX�:����������a�c�yS�'N�h\��I{�gį�4����ȡ��kϯ����!����/��J& l�j��X7�N�������1�d��z� ��7�B�G ʔ�Vg�U@��)Ɣ�0A�r��T/2������x޹�p���D��l�@��9�ro[��x�5
�?���/x������he�]Ke�L ����'�Q<�,�A"w�幉L:�} �a�k�DcϷA�*���og�[�nNph�4}Ѩ��x����5h{��e�=/�tԃ��ǣ@����#�f{a���\����G�l����_*�p��
��ì��P��)2*J�D�	�A�MZHn�k̨[�T�gL�șTC�iS��AL��/�j��6�3�82b�.�\������)[��I<6�<ʚq'��[�F��
)�
"������E��rx�~���&�%]�=��M�,� C��a�'΂#��=P�_��d1'�/�$,F�͚������ĳ�0g^r�+�	�KRI���)�	a�=���|.�S��d���r-�8�qv���E�~W�TQ��ޫ�s�៨|��N`���:7��IK�J�]e�����/��#]���Ԑcpѩ��74M`�b]n�,*T�Z��XlxVHYEB    fa00    10b0���l�i�2�ɰ�},�扩��Z
�F�`1A�����6�=���l�����5�c�)��m��~��܌L$P�s�&��QY �``�JE�A�[8����F�6�X�>������Y��n!��b��S~��y��"^49�f'�	*��0��A%n#�B���q��ԞC����6��!������,�����~M����7l镏<��nď�6d�~�g��`}\���$I|�*���zu���ϐe������M���w9�=�3�F��*�z�����]�+���~@�b�v9� �/A�4e��)�Kp���vY�����04�ś���N�,*g�R��5S>Ds/f��ŕ&�y��+�O��P��U��m��W쳊p�kh�6%M��^�X�vM/�i�+�"�_:-�� cʒ|�4�9��;��W�ΘmD�轘��&��(�҉�kº�R�D����8C+�ܧ���nq�=@V�{F����pDr3�1?S�c5�O�+B]@���#�*�ׇF��g0�r�S��^AC�(��H�W���J�L�g�-��D?���$ſ���~�Y�x�?K�s��n���)7��uW��Ҡ��@�=ǘ�'�]��Cf� ����`v>�v5����#'��������}z�ٖ���r5���jK
7_cճუ
s@�� \"%����οNz��%��.�b���^�5d����?� b��Y��1 Z�#识$t��3�#�ո������J�-��ET�]����Ӡ�0%Wa��"��Dqۤ|�'����QWb�����m�[���ch���Z'�Iu���s�?�i��5�bR��rhD��y������Z�;y���5�q{j�f�m2Ĉ���Ebli1i}�}�FTX�ր'O`iաyf��m��u�Q�u?p�n��mn0.�1�=Q����f0_��}[-F�㍋���#	y�� q.��m!:���:�h#>6�vʶ�s���C �+i�'�.s�f	p8�W�_�|^�%vm�жH��^&�%��X~E���u�􀈫%�S�[�6߰^��щ1�چ�JJ�7��"皘n�+��>�z�q�/V��
e���7� d����n��*��?&�#���}|g�'_S�:W�s~�9��^=d�Ev���0[Ǆ�y����Ę- (%b)Ұ��dvBX��ec,�F�\����m5�>L�IY���_;�r�}�U�I*�;���!ߞ�o�ːFv������-a	��^��t���� Ϟ�l�t>%��cDj���҉��XG��1�7�YA����H��>�{h1!���?Vȗ��'HŬE�<! ��,o�#=�i(��S�lzЗ���ԯ���?=O\��� �m�X��
�~J�v!�������O���VH����R����*�ތ��5\��&�p�~��'��;h1�5���E�J��4�_��"�p Gd� R��"�ӣT��P&���i�T��XG
	K��3���J/ú��;4뿾Dn���r�-�>ط�)����#Tl�� ���K&�7 ��]
��O��z�wj�1GL�rLU��ݟ�A�J�����m�È� �m)�[o�V���aV�B�o{�D���%F��{�4�� ���*u�&�|ˀ�_B��+[��$�_��h��{�B���a����R�ܼ������-z�Zt����<��N4@�,�#cFfƯ��@}�*�L��ܥ[y)�I�_�ЭM#�#~y2�y��en���ԱU ���@��v��.1ܫD��2U�9:�Z�����4���Tt���ȫ7:4<1\�9�zf�SZ\��~D~gY�������疨`xj���v��л�n �/���Ʃ���h���r�)���3W ݚ�%|�V��`ʭ����QLb�ع��ξ�u^�Y�T�'aO_�n�#�ޠʠo��AnȢ�Z&X�31`���c�--���0�Gq��nՋ߸�'�]2�MO���u�����3}�����}�P��V��Cb%��"��^�%l��X42l�=F�Hm�s�8��g����]���#��O�Z�ꢽ{x,{lr�I�a�3v^�C>%��,�����`�Z�Yp �06���pz{ωBѭ	����G�Lr��F�*��Ck+N����|�r�x�в�$!'D�G�a�wG����.�@��������)byoz�:��f�Jh޶�ҦѶ����Ӵ��g	Y�����9��G�R��{�M��ʳkȥ���P�������1����ֈ)�+	lJ� �-ȱ�Cc{xb��lͪ2Z}z�Uh`�3����6rCV\��peIҼ���RS��B����{��:6љm�_��o�ګL�'j�|El{*�n�V�s�o����5Cz5�N��3"��-R#8L��`Vmu���|aY*�
Vx:�~�Q��x��5�h*#
|s���2����'�<�k�L��nUV%�3=Z̙/��w֦w�*y�|c6���Rv��5\�鹤_K�J������0�T�Sd	�1L࢝�78��ٮ���)�6��S[����RY�\ŕ�Fx�TF����\��#���M+�����)�*P�|���2?��d� �}$���h�j�b(�WX�B4���(,�9��y�����y�!�-8�UrX}�!2�b�;fX:�C�";��G�.�Y����6����P�:���]�'�*�M���
�~��IfS�M�c4.%jI澙
k�͢���綽+���ݭK�o��OoUbg��N��7����3�y�#���< ?��v+�/=��$BQ(�]�TFZ\"E�^����[_Kv�F3�����FU�ꨌ�R�ߢ��t��bf������Q�dl^�� �o	�>�N�0Hc/}�>�
$��޴�B�QC��œïe)&�uD�G���nH�[$diT�W�R�|��o��,��68���^?�������`?��x�Q��U�cC�P�,�t�� ����ui�ty�|t�
��� /:c�-�ۉ�X�Z�2��� }�1�ZD�nͳa��#�T��O� �����m��"0_�$��p��A�;(+�s���|(��ٰZUhk�*�[ffE}�!;���dcѮz�3�z��#Jw���8�*?��k)k�(��󫯂�[Z
oQ�3���w4�e��w�O�t�GlJZN���Q臘���JKj����T����k�<�
'ʆ�罠��F�sɭZ�R(Mb.�'d��ՉU��`����{)|�b�9���0��^����{ZW�w6{h���O)|%�l����M+)S�?�.�3���m.6UW��S��g�+Q�1��<����>�:� #;xp�^AZC0��ꞇ�LPwퟌ�G%.�|�!�N��mNa:M@�mfxSBNA�Yw��>��㰭E3�ur�PE�WxPS�)��R�`o�gލ���"�7�H��4��Gz��א)&h. ��1�<���$���F�}qW����޻z|W&~�(��d�C�P%]Ax�a����?Fv�Zr�WJ$p�V$~g�s���/�]-�S�pAPG��M��Ț<s�a��Cr���/�ɖ���n��1h;0K�80y|Hϕ<5��,iL|no�<m��KN�uQ�&]���7���&��[W,��x� ߫9�����>���l���DQ��gIDִ���X�۟� H�=_�p�Tc6Ry��4'�(�{Yc!PmL'��S�!���	�of!+��z� �t��uب�:�y���L�,�@��_N����]���o��o@�G��|��v�| *L}����Y�~&�����.y��F��8oi�Q�qፗ�Z�k�M��f	��A�܎�Y<�O��'5��3�́��!T��'�]R��S��n*
c�! Y���__�%�>��bSDO����yq��f��Vv �8���dE���	��8�]�f
W���Xԣ]N�Y��]� ��,�S�/����ϪJ-4�J�V�eb�j��v$��Q�=L�<�;�G�����􁮖����|����"E���6��G��F�����9U匩h�@'��ͱ��}&�����bG�DV7��P_��ѩLq��nA�Ҕ,�x�k�:�?�������M�n$��՘��G~\�aJ����Z�S�P�K������xɤ�'�Ć��͓/m�fe��O>�&ʮe��C�b▙	7-���,���F�XlxVHYEB    73ce     760�I��t���Y-k��#��ï����ld�x��In^�Lu�-�0m�a}T2^��t�-�ݠ����zaX�z�fN�p���lPE��
L3|!���r��nX1�`_Ed�V�lP(q�G�筕1��֧P#��kzz��ة1��Os��e��>t���~N0�.�I��"$"�Ӥ����f#Q
uJ��~����; 0��ţ�oc�"�XG.Zgj�8M�� ��my68����H���������{��KU�G��$�kW ~�lO�E<V��7+�IV�0E�:�ۚ��h惁�=L�OZ3�b���h_�>����ʊ�b���s����n��ֵƍ��&U9�L7`ۦ�W�c��NfEΑTF+�A�>]��~�6�j��ے@)A��܀6M���9���#g�2�D��<�j�,(�
ô�]�̔(aEt�$�	9MlrV����]@!e��G����K*�f����צ���}�M(�ס���D�5���j�>���i�i�.�����NM>t��e�pzS�N�) @ge��Yr�[�A�Gus[X:sڼ�Rqo�ܨO!�5�"-�>H���ʌ�	�pYI�/fP𓯚k���t��s^w���ځ�����Y)�Vl	�]Ak���'.�����4�_�S�/��K�9ن�����󪷩�F�$�vbNi��{��c!�����c>*s��*�
�F��s�#�O�)Gΰ�e�9��3��`�3���uS��	 @~�c���.F�g�O���f�R������IA3x�S6�{�p}���TD����>��6$�M��/	�u�biiA��{�f�8`\���[��DĈܾ�("��;��k'C�)m?!�~S/��X��"��a�U[#��z���� =��%e̝�xQ�yH��ê{�*�i��ch0,�
C	�B�:B\���Ϭ�q�TS�����NO�>}���T&��2���1]Y5��{��gi�� ��C��C�pK?(��a5��=�ԭ/(㕰	���ɷM��&�7��"Psw� e�	��3�	�~c�]C,V%-�V�sf��	�_ �b�G�2����\/�6�r~y�T�	��2�f]l�k3�8n��p��`!,qͻ<U+-\.Ȍ��>�j6�l(/��g_NF�8��7ns�|�t�m���������+�.!Si�썒o��c�6CA�!˜��æ7F���<��&��Ľ"���c|*�r`[R�d?�ߦv�#|���wC����Pg-1����R��BFK�7R9#��-J��(e����H��{*׆�y!�f��ɍ#q�i�/�CUu���Rj/fW���w�i9���v@���� )c�ƿtӑR�����+%M��]����Z"�`m����`
C�.v �g��-����R�2$��'���X�C2�q��C���/z�W�&W��6���B��jcD))\����d�����f�^❇)NZ���XH��R4��+W���LX���7��w���L�e�O�����4��Xo6P�{�@H(�l`>�L�h7=Pؓcrk�q� �C�<���?��ީFr|��kQp�.��i1��Ū�8M�GG��ͬ��^�hR/�L��i�<�n�o�t΍�(r�*�~g��d�1�n�X��$��l�&�7�H�����Q�g"��`�u�����Ӳ͓�m&.G'�l�,TB���r�$Q}���p�|X��n׹�$�{���5�9JY��D9���Jn* �'�
�Sܠb-�%���Y�����:(6��E��],d����~ہ�ܫ�J�X�`��q�gE^�/���������m�"���Mէ�V�Iܚ㪵\