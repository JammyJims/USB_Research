XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p�iSS��z�*��z��Js8&J��#1v%����#on��R]Pg��*0+���Q-$�*�j*p9?�;�ㇱ����@��7$�魙O�~%_d���6��T���1 ���v�C��է_�p��;�0U�������j��:��NҢ?W�  �u���#�g�0��(�=�� ~Ț����-&~�,�g���C�~��
�CeVǑ�����X}x�!�ˉ�P��i��k�ر��Uq��t�7����c�P�K$�2��x�0��	O.�@߯�S�ljcj���&̈������e��0σZg8z9_('��n�[j4Y<����E E�+_2�,���G��B��� a���/^���R��2�����{k�H��4����D��hK�B<����+���D&Y]N�>~ZR��r�o):�'��X��QKrJP��$*�B��I����*�����GZ���Ot�b�j���=�a�a�EB��9a�	[��#ʷ�*m��\����b��N�i�8�L}�׮���#{�!K�m �2�KY �F|�B�wh6%��VE�X3<U�r6��4��2Kǀ��+W���U
V�on�,��J�Y�,�ѝ^^l�d8�<�]J���<�a��t�	D�őf�l����-��� �s�T�#����5��6P16¥�°rL�x�K/γC��E
lN�5���28v'`���#\�霸�-��e_c)�I�>{xcVO�.�@�F�RUɊsy�e�XlxVHYEB    859f    18f0B��oa�������i��?��[0̳����o���
�9i��!XO��3�C���$d��[NlґӢP��_�����dĩ
֌��3J)*��!d��+VY��Ѓ�q���|��z��wc'hZ����4�A�,��f��p�>y-�7�KdI��<���Vt�� P-���goY��Lٗ�|��Q�1}���7k��7���R#�W\���M�	�N��ʈ�%l�9�Kс<=2`#��Ԯ���*�(2�E߁��,����"����S��~�%�\d@P$_��
��2��pm\,�Ǚ@dy�M;>XاbMB=��[�ƿP�&��Z[#r�vS���f�-b��y����
b�k�]�9x��:�Q�tWq�NC'�@�l��mYe"��l�*%Wq��gܾ�d�e�9HI�%@��g�-ɾ��
�&%�F*	u	��O�G�Ʃ���I����dO3	�?����B����ܯ�dh�b`���������E��|r|���)�%f�
��2�Ƙ�b'p��+�9Z�/D�bg����~��QyB�=�����ÿ<0:h����o9H�)y�{2t�Ю��Ȼ�[��ѽ��Qۀ.j'�"\�Gv?\���i^�.R��?gm�v�RV�����'�x�HpI1=�v���)⹱D���挻�V1�\�8����%���^�.��x+��Y���y[
j��BW�v�ɖ��gJXG*!��������+����	��p� ;��,un�ccH�Sr߈�,H����-Y|���:�����C�y�_�pD������APNdg\��R&�/�EL~��G�vFk��Kw��ꪪ�~�e��xj2����������a����/�R�x�4i�4Ќ}��2�/�)Ѥ��z���_�`?��6�5�$u3U���RA
g��IW#��co�J����[���^�|���:��!;i�A3� 7�K])�o���a�~��9x�.�6�W�WW�����]�ַ����:��i�++���'�F��Fc_cv�$:s4Z�Y8e�q�q�s�b�r%iWЎ���������sЮBK��x0Q�s^g�ji:�*Ŗy���ą�b��:�3��C!Dd��4������<ھ���
��G�!f=%I���:�Jv2�y�d�"d������ߕG( Vhk]��0XC��p�r�?��J;�����n��ON�hJoW�4�o�@=��� �V�p�x��L}>�_ת��0wBb�i<¿�SU؆����nQ��֖��6|��P��]@�Ą@�߮��=Y�hs�<?jK$�y�Ī�?���y ��8�ă�����}�Y ѻzY����i�<�Y�/s�U?z1����ZZ��T\�($
�;�0S�b�o�0�q�r��̵�o��%2)��1	˴��Ō���4���EN���ߧ� �-:CZ��zgi��#���m���8Q�:^��^��l����o�%�e�i�_�M��[�t�(��)���D#�	�]���S9���f�Cy��g�X�߱��Efn�i��L)E�-=6���ƻӯƷ���� �I�bYݷ$����Li��U-������Y��xW�Vxn���8ǯl��RR��	=�,�Ty%�%~k!mЏ=�S|��A/�a���k{�S��K��Ѓ�m�#.�}w����۠V�<�n�G�R��/:-��GD�{Xش%�qbu&����`��H����dOݰ�&��O��6N�Em5|��ll�,�������̈F��?$�h�:,�o�rtb�PP���ڔ��t��d�i��Dhn>��b'�r��75�K�#�����eV�ʛJ`�jN����rHAfي�|\m�Lا�h�����E?g�p�T*���m�͛�]���00�,dF����1�"SX[�[6��G 7��yp�(�@ģnsV�%k�hF�9N^���&�M.��:����^���Tm<��|D���8NeF�:k:_���Q�yݾ����N������p*���PY���o2����.�����\>�d��?������m��F�A�����e+����n�]8�߯ �;�$>z�,�B+��c^@�߃��l��ެs�}��}�SN��耟�D�篠��8�%�5��6$EMa���;�����(��u�H1��0��ۃ<K��� �Bv/�]��;���5�|b�P���gfϢs���S�}���&�ֺ�
�a�M��t��o#�`�a��%�O�ʢ�6i>�^�6���*T�V�)�YA��c���C�a�� ��O�y$ߋU�ϣ�����J�3��s|�u7!H�ـ���YC^�4�"�!�b�i�(�-
�͔:xĤ��d�� ��gI���KÊ����ּ�����^���L��,!;� �:�R��ԉ'	����b������l�7��YPz�%v����7��s��m&�qZ*G�
+�H�q���% U�D��j�Ĥs�rǏ�����YS�#��Ra3<R��r��>p'<�o˙}Ⱥ�®�h
����m��i�e�?�US���egw@��Z|PBM���a~����m�'.s��}YJ��kj��p-���t�V�1%|V���@��#�!�}ʁP���5�v	cm�D>�w��G��8���}��9��nG(	H=G�XƇ��A�
]]%�QM�Lh��C�����F����v��Ώ��^�����tr����CGȨ��:�.�l��`#,Ԅj�bSnL�*�.z�4��zp� �2*бX/[R��؃"Ʉ�f�׍�� ^�e$��(�_	�T�;9��߷����l��������]C���B.E(M�zz�0=�ࠋ;w��1��MM�j'Z��Y�`D��PY~S�V#ĝ0K;'��o��� ^��%�몸��Ly+$��aޗ|�B�w�w�ٟ��"��~k�A�ˋvˈ�A�ן��Q���'��g���7u��_�7=�����;���'u^��9���R�٭#*�"`,�'��~��Tm<����PE���PL�E�����ѾE���HK)��ι#���
�R����+f�?��'���h�Y����EP�?u����l���z��J5cm�!w������u�xaK���ĞC�@�i
]����z�{� �D[��j�6E��W��{u����Y�Ӫ����9Q���ҟP�� �y�z'|(v�!�
���\���z��/c��	x�'���3�$
4�F��!��������Wf-���&�}�yW���1���>Q����[�����n� z�R�+#&���X�.|��so`yl�a�;u#(�ꆄB�{$d�C9���Z��q���~<=rk>9�3�>ӎBP,��d|�;)T\n�J/	S��;sQ ����m4Wzݷ���"��s̶GՂf�t��ɇ�T}��I�)��ҏcSK�]�j��w�a��wp����`��nNg�ݒg >l��j�)�V��$� �d� ���w\3X�����y�S�g̡/7�������G���=�=N�2�&��n����sP�_��7��%I��I:m@Jh���v �R뇼)�r�t}��Iϔ��ڱ���'BR ����*3�O  � s��E�::�1y�-Z�]��-o��(�r�qA;Ъ��HK�&�;�E��|��r(w�F#go9*���c�ƥvI��،�"�ؙ"�f'l��P�ZA����� ݵ��UH�K�k�����D#�eU+'l�u�=d�5���[�_/
b�^����0�y Z�B�q #*]�8�] �'NoA�7Ax��<Wx��_!����C�O�߳��k�i�Iw�Q�$��`l�RY�4�W�����2�si��Ib$����W;�4C�j}[Y~����HaeMrV�����y���Cod��C`M�n�~~�tF�&(Ig��&y#&Z�c{Q?U����,IJO�[�i�|�dGu�y)�Y�k�2���9��kf4��$H:k�H�)z�FvoQ"��'�4��1��Ě'�lC=w���ݒ��L�k�'�[��I�{�j�In̻En������H�b�hxzf ��]��*�����~Н�pb8p�f6�iط#z5]L�(�$�z1�f�e��M%mM��-�Ӥ|#_ŋ��?��5����EP�I����zX(���֠����*�DgK���e�t�jQ�[��,G��Uq'̈K�E/5,8�!�2i��گ�s�_�ހ�^]����S�i�f�i��'J�\��PZ�Ʌ�p�Q�*�~�[ݡ�mie�l% ��������^�:V��l����A�����)�� ��R��O�]'$���0� k�v����FmQL�r��oX��9$w�^�&�9*�@6��-���+إ=�A��̎#����O�ЦObx����O��1��
�nu2��"6���O`�)��!6W�K�=Q�a��m�j��7�i
�8fx	!~T0��t�8A�a�6|�����6����<�G˚���a��B��۳��!�mj�moTr���/k������D�87����z>S�oHiWc䒑HCgSq2��>�����������U�F-[�T����u\����N�!���Ԣs����������(tvz�|�E k�/�z��n�T���Q��L�G÷�J&�~����� @�_�"!�vF�";�J��ib,t�=ȁ�����38����Z1xҊ"�q�����+6�b���N��یJ�23 ���pPk���Xۜ��S����gYS 1N����(M������`����	����S�B@��j[��갼)�G��3��8�c)��?�&�Y�v�rX�l�@E,\�B��;��=���Hg�L\X7�����/�8�7� ~���5�^0�����c�����hˇ�.�R�T���w۱(m�i���	�@�a|��U}e1�"��n�UTh�p�һ54`���^O�Xg=|����cf��)mb�D�0���ڬ��P�4\�RҥtN4��q��8��oWm_&+��x�_��M��`sY7oSz ��h�J���0��v���~�RT�'����T|��e�Q8c����	���l�-�e�v�&Y�VxG�̳�̓���pf��\o����M�Y����H�,(�!V]?�����2�g�'hh��,{�5�����o�0w�F�x˂��.ѣ���?X�v�'�
}�P��3ue��'�z$�,:}"���1.��R8K.N�R����Ԃ��^��B$ <b4�ՠ�{h�ɪ^�rJC���-��٫���:�W*4l4�n�v�pҖ�W~�T��JTژ��@�S���G�jT0��H[���.R���R�H����|U���M/1�Цi�]:�A���Y"�%�̲ɐpp<p�F���▏ܹ���t5M���ʞ����D���-N�O��#�'n�j���0ss!9^��)=�|p�����ȃ��d�;�����4O���H���m&�G!��B�6�ҙDӟ���,�C����s����YR��~�Ht�|5{�4wjr��F�𲣈|{�����@7��;^'k�tASN�Kt�L�R�m3��i�է��3���4�M�.��+6DS�?L��1����@-��g�{>Wc��$����)B�zO�
]8��#���6B9W%P�	Z���������ִq;Gm��C��p�V�2�|�l������	[/n0�� �y> ���闡���$T-����L{Q�)_�z�l4?n`��c��쑵�b�~<��}b�E�۳2F_�<4�
�r6��w`�;ƨ����^^��Le�a)�����|<��q�[��P�ؤ�~��Ӻ2ucY��C+�
9�iC��Gc�G�]���c����o~1Hr#}��ӈwUw��1�O�ܚ3c�>OR���]�\Q ����8D_Z^��=o!+\��.�sْ��̐ЙX(#��`�WG��%Gh���A��+��}%*�<+حk_y��F
$�:�hn.���܇-p�G9M��i��_H�[�rI�ج��L\�H�P�g8VϚm�Зs)�S�ܖ8���F��۹���W]t��\/T0"��v��qq�YA�d��mϼ�>�HD)�G�}�2'ţJ��P�c�)�׈6"�+3����њ�M�����U�7���T�.���r�.F�RAI��NF��*�xa�m��6hw���O e����Ry.,���ʵ�6�� {�u	���zP�p٧�m�`p1˪�=��T �^��0�CZ�\���AR�L���=m}��q�Kp��>�
