XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�V�|�Jm��p>�<pz�1�U�t�K�$h��j��uK���cQ�3���z)Jj�;w�@����m��.�4n/�܊�P�gjO;A��Rr*��%}�6��U
��.:��Z�H(��O�m�-n��D������Eq5}u���tq�!/FD��ӭ��t�Q4��6��'Æ���O��(��ND����� �欬[���{���M���Io1![�xo�^��b.����xm��K�-��9�� @K��NÍ��[QG:�c�e�w/(����jCiy������I/Z��+JT;z-�>�K����B�N߰6��=��"���sy( �X�i��P~l��w�;ɜ�[˟.n��3�q�S��F��-�TÁ�7����Y�}������j�\��e�������0�%f��*��a��� zp���3@= �����"�Ir�)�N�L�⎌�Gϣ��F��n������+鼼Ns����]Z�|e�����6i5ĦA�Um?�V)Ox+³=�Ny�2�%`�N{L޲�KK�7�3��|<|�5x��n�����,��s���=�h
��&�[W5�v���O�2H���C��f
���Ѫ���#���]-��YE��	̍�m_����4~�PG���=V���v�r�����-�"��f���|�X�t��S{S|�>�i���5����3P�d�f�"��N��8����.��;*�:7�_�h���aa� �'le%IT��h�BGC [��XlxVHYEB    3c04    11102�:0��ɱ����#@�b_<&��ڬ����ьew@�>���iD�og��c�t�����xe�nDUM=N��g�Z�T]ڕ:W\d��r�Dp5-���N�e#/��;9�C=�(��I�&��=�0���~��2.�l��[Tn~k9A�_%����Yx��[r9�M����#ޅ΅��%�$�)�?)��<�ͧ=�dt'Qj^x��̨�*$I"�GJ�"���|��Er)uS�'�{�<��Yi|E�F��x��IN8qۅA���x*s���
��z��q��Wa0���g�@�� ͍����G-����ݯz�$9@�Q��{ؙe����M��#1���� hO%e<�<H���7@"W9+z
��8ZL�u����l�j�~���U�,�����0CH�յz�DkmB`5�����e��>6q��/Y;��gdb�ѧ\CL��=�~�+܅���'.�k�9Ht޵(�8S�zqM'�����82C��L���>`���+23��lg�Jn^jʠ\�HS�|��Y�Cj��Ƴ!�M!P��E��f���zگ��X�J�>=,hʌ!'[��:yS!Q9�)ʎ��r�*�Ĥ2�M�O���\V�Ǥ�"F���2��lFU~uD�Ga-"��b^Alnj|���|�G�o���������X�d!�|���k����aSpV����?�w9V��p ��{��.��=z'qE����x�$&~���<_s~���i�ÍE^�x�k�Y�j�6��%
\���\v=y�ʎ��}�y��قl�����y:��j�A����]+D}m�����S�Lj��K�p�9�XI�À�B>�WF��m�LF�q��I8���+�@�p>��R���3z���3�3�0�� ����w��qsJf����a�#oշ������Zۗ�pw�԰D��p�+G��[n�  �A|�\�&��LP�c�, ���a�����v?�׎�U��HÒ�0���B�gR�E㮁�$�ړ`�D�tjE��n�U�t]r��t?q:e�^�3T\-M�dYv�y�#�����;���aM�8�@��i���_�:�M���u���2c��ď<��� _W��v0�{
�SDhƵF��R�Kݶ;��$��Q1;\�]�4����M\����{G���Z{W
�<��k�e��HUH$��L��םP���}ǿ�4f:�)���2T�|���-��ۙ�ڑDL�|�W��ܳEe��M������b��E8���X�`�v�)V�Y�������Z_i2�GYc�+�D��ڤ�l{ZlϯI��̫�G6���m'�ķP�����=!�+7�0�ib.�}������vG���}�<�4��9��文Pm�o��+�+��p�'@��3�b"*Ϛ�D�F}ֿ���/����B�\5?����iC���~��~T�(���D�DiN��.�`uO0�Y���4Ç(�MFK�*o��j\��f3�8��0�d��a�=93Df1Ŀ2��o�T1W���o�<����)�-��[H<^R��������24{���.B�x]i��T�Q#ʵ���)4Dk=�J����4`����-~��Ъgs.8` 0��l�3�Իq3�&�����=��M+d8� {�֥!��Y���ekj-���k�yUSi˙|�p��L��G/�� ��I��� '�d��It�9��.�*P6u�C���Y���j`8X�]!�[�h�D?�L�^;���2Hͳ*��t�Vu!��ː��v9%RZlx��S?m���	��T��Wt�8<�`4�c�,�0jdm��j���c
�J�RwlOz&vɐ�k/u�V"jޛ�x��:���N!k|���)���~[Hw�4���`�5,UGo��}3D��aԴ��w�]�CvP�P��.(O�l�.0!?4�m�U���dC2!���%�!�����CeX5*�R^mo�������ݫ�oy�uk2}c	��vA�A��˫H�� �E�	m]�W�P4H�D�[1\���M�/`|M���/�����Q��5�׍�'�;��9t��|x�DP�`c��2n�toܛ{{�ӹh�ݒ�l��Hp_K�= �W�_[.�P:�5�T[�{�͘���=�9!RY(��R��)�F�$*���(ˑ�e,>��*¥�A��˾5�Y�y�~�����J��xĲ
g�����PY�ĊSћ�D.��!���@�KLؿ>��s3pٶ�J� .�p��A�pg6&7bVi���Z.5
��*K�1��X��x;k��:�y]��0��̉���6�qv�������L��9'�(���}]���6}�Dܲ����YA���;4��0�w����H���[����c9e[��4�-Y��_��"�I��������5ĕ�O�E�H�1L�#Z�s:'�D^8�=��5���1j�
kJz���rs�$�K�F��w=<Ky%�u�Z@xK�ۼ�/���djt���E��i�`@s�d��ƣ��i0FmX
�)iĆP�G�
\&�(�@4ʞ���Z�/�03����[��r���%�=}p	�y����yU�5�Κw
�h���|7s�Ք�R���g$uSr����0s?w�Y`��ƚΛ����(7��&�┯Gt�O��B����鴂�y�CU5f��_%ۛ���gi�"���'��/��+K�����{V���������h�D0x1�	d��<i�3���tں]-� Íq�\��%n��:�{08nM�J�����i7s>�&�((Ѿ9����M%?�~��Q6�G:B�pW���+�ٸx���Ri`��<�HT|�݊c҉��(����� !���
E�ꏑoAOut��K��nLERTHFd=e�8!����+ֽ��ͣ&�*��}��x*CFM:����?h�\�2y9��������$=�ۼ�~�,��t�H�����o�#��/eĽ&��XQ��>���? �7�7J�;t�k#�Z�	#�m��M��F����"��X
co.McsR����(
h�3���ִ�G�4���Q1w�j��Q
�T ����z�_�����OՌ#|��?���I�"?�2��R������\������3��J�+Q���5�Te�Kg�r;���0Z�|I��g��M��=�D ������m ΁e�Ko����~�1S�O�t��cN��@���-�h���)"�rl/�e5+JPm��r�(��LɄR:�>�ێ�N�|A>x�j�+	,���_��~� ���_W������'�]�b�.?�.�3�S��ï��q:At�#P��1�{U�.\3�N�vŽ��UMx
*ρesn+�Sml1ܙ���R`ȓd�e��j%�!�g��2k3&�W�,�>�3 ��a��U"�,R?YČ���_<�^����D<Zۺŋ�;'b'��*lވ�E���u�Ɖ��|N������^wS��+2x{A�R:� Fڎw��3k�-��������3 P{ׂ&���N�!*@�-��P�o\���r����Nj�Y�I8M�Sm���[Nl詊P�O��%aQ�տ���o���!�C>iʁh7���jm��"��<�|W3�('���a���N�K�a0�p�]���Eح\�)�
�9�����6��x|owfϛm��O3��;��F��i�"*N�6[�����a��q;+�a%�r(��PO�އI	�b���i������tG%������؋�R�L#�5�m-�\N"��LlJZ��pF�?('>���k�"%�e�o&�~���'Mڦc�I�h����R��^��2�u���z'�U*��D[���W^2k���0��_9퉱����E:Z�z�����������OB���]FKf�b~йv���R<I	e�|#���:���P��)Z��D�	CfHN�Қ��a���e�\6�F�
��>m�e�I7�<�nɬ=�+Hg��n�2��q��F-����[�Q�E�d�NW���pE��yjHO�K����3)0=��,٥����Йa���(��;9�K�P*:��w��]�\4�z�~��������1%3
%�:�+Ҍ<I�pg����x��w�D�2�k��&]iEf?���V� r��u��1t�>Pe[�a���u�d� ���2]3<��E�Yᛎ�����D�"���Ӎ�D"���ے���h���&�*N�%�A�Dv�^J!��y�`k��h�`Rnя0E�4^���rr���u��0�<��%�L%�%̠��~��tz&�@�"I�(�g?O�"f��Le;�\3��]��QO^s	5o���;�8:��K"q)&�2��x�b��#Ե_u�0��