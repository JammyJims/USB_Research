XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ԕ�˙t,�}�u�~�G�I���O]��Q��he��JQ��F��m^�__ƙ��ĵ�zz���S���o�a#�\yh�̪�����j�R�Ԥ8�z;?18����5���^�"�����r8Ҡ��v{4�aB��&�I�H$���l?��z.�5���@��o����^MN[MJ��N��	F�í�3y�R/�o`�?0�~�j_[岑I�ӊM8��5=o�u��̽�eДO�	�,���c������X� �E_3]�$��ˀJ�	��ݘ](�D!�]D5�������f�[�����KA;���;&5�?Boٍ�k7f�&�r�>�E�Ai�j8��R�Fv:1��T:�WOPc��[:�I�T�V2�.���e���|��h߬ۏ;}tvLijU'��#�{���n�	b�3,g� 8$-E���M}"xƍV����A�t���O5�i��,
k���5p(=e(B٥g��/��Q�Z��d���������1YY�e�s��7$Z�cf�4K����5���Ƽ�RM�+��{�⩖�s�|�GL�y<ht�}�B�)$}%ɧv~�����[�u�B�ؕ^�g4����C~��:a�XɅu���D����$̛�\�F�[f/���N�ˣ����+�"�G�
c^0���\��@��?#��]���v���x��i��v��h# {���J�"��R ߻=�H�Dϟn��6���+-F�TXlxVHYEB    25cd     c30���$			j��p}%���&I>U.��Kf{4��64�`cФ��W�J%�b܈��EW/}������s[����﴾�	�QTO��D3�}��������~C��6�Pn&�@��F"}�\�̞�|�<� ���@�	�qHyR]#�␇�W'L����A�|TBŋY":�-=`�oO�m)��`�qFn�� U=�����q��6t��t?u�	���_��DoY��!R���j,Cf㖱��*�b����}#��D�����m���p|z3��9m���]�&{ܴ��:ېb �*D��֐)i:��&W����{G���b���L��F����m�#���1^b�/�j7!!��b�#Je��g��M�ވ/��Fǚ�����]��D�������|@{c�o�$������ֺ�QĪ�oÌrw��i3�[)&���?�z�-s/&����P�l�hiF�%�L�Q��������y�p �b<U��ݬ�/�@,vl���wG��,Գ1nF98����,¬+J��Z����3I�pm�y̅%��N�ߎ��+C�c"���6���=r��ַ����0�`�Jxϋ�ǉ���X��#�}�И��݂�Z����b~F�|B�J`Dx��T���;8.��'Jt~1C[���ȸ�~d�+�	6�:�b
#��D��D�"�*�qY>���'7MH�T�\��ګs�l��>�u�F)�T��̴�����TO��8���$�T����LT�wxDA׉�q�A��j��-j�eh%�!�ݔ�z�����W���\��l\J����w�����+s����^g<�W�=sB/����?��4JV�Nު�^��c����I�<<���M�˱��54�k0��Ɍ���@mΞ71�Se�f)ͬ�m4��J�	�.�_�vf��p�o���}�VEF�T6�28�$����{�ѹ��$҃Ñ�}� 8�[8�
���eX (�����y��+��KV�`�$��k���bW(�ҠkQ��xP�D������Ȉ0k�E�u�p���S�άPX����&g`���P���cn-�Ǳ�$��w���9k��f��o����s����Ô��	��Z������p�gw�w� �)G�2F�Ph�+��W:94�_�o�)���2���[�ʮ������˵��	X�h� >Ao�#�/Uu�?�2a3O]��j%χt�ARr���P�ꍯv�.J+���*[����Vwɨ��T=7r!^���nk')񙦖����O3�a�MVuÒD��w�:k������Ѕ�{�~erD�i@�`ݕB= �#>J�T�x8�3����[S�7b�|am��Jg�D$ًz�g�/�WYf���
&�ʯ�����u�ؘ�"���rKƯ���.I$c})?�"P���馀�Aj+(����	�D�4��AR��GP�M�O�X�ʙ2��T[^� G¦�)(���:����J�N�ȧ�.:����_��� ��C�O�����Bg@y��8��w��D�Ɛ3r�����{���e��PP7{;|S] �һ���m��q�GnG�����<	
X������؍�Y7�o
�7qr��9�#��p�������F_��,���Սk
��Q����H=�8�Ӱ���)�E.��Lq��J�j��Ø���n���64rVѯ:�B1�*9��,KZ��)�[T7u�H](	�:�種��&:@j	��K����Jt�v�/�Aaȉ�5��*�$�\l
�g��<2�>i}?��������[漖/Ў.ͼ0`$�R�s[f���|�b���1�_hrOp���+ʁ��S0��K��'�f9�:3r�m����_����FE͟6�[�����YR��V6�.��d?ZST= 
�Kh�߅�����ʰCU��!Ug֞6��
�&Q�2�/|,5KJ]��t����>�'�L����]�/���\��>c�8�o�{2�����} �1����\]�+�(B� ��P��9�I���G���b�i�e/�]��J"Ѡk�ĲL�Y�n�S{:�`a�����ܹ�o�8�P�>�'��/P��ʌ%j�*B�����I5G�ֿiX���[�Pb����V�by��^�eMw9��J<6�@��������;����s���%e�
ܿ1P��4+ �D�o�Z�Ҥ&G9�B��W�"�9+uI�蠯A.�Qg\�,��b�CM�*��(�I�̰�Ζ�KI�}��,L)�:|f��ȝ`'�ͭnT� pi�H���^7��Ӂ�#ڀO�����=������k�F�Va��)Y��!��l�莦�$m����3���̂�!i��;V�!��������K��ES��/�4Eh�aFG�Uh�P!��r�ڽ:tCW�wh�x���X�`�Ͳ���J8N�wMAT��PIGD���
�)!脀��= �lE�;�tBLXz�i��}�6M>�/.��1�񃟻K��,p�м�I>f�I�_DnR�t�,6�W�:��g��]�n3�kI�7Z�ꁥw�V	y<��8&���WKl�*�r�xv���R�~����CAd\�O�:`������� �J�9X�F��P�8�f�k�T��Aw�vN
���e���N��1�=��3�1�b�1�r�F���j�Z.��G��mS�NP���S[�fA�g��l���g�Uup�h��E�~]" <K�boR���I�/w \X���l�B���$�K����)�kIت}{/1a�l�7Y�#��Gv���@Q��:�(W&�p��|g� U���2��v,��f�n�B�3^�O���5����6�Ľ�c�x\:
��n��,;���z�e�M�:�s�n5�%�8��"m�r���Zp���'pc�5�ƺ���/]`�SwIP��2FL�=t	��ޝ�R�f�*��-Py�-9�G4�<�n�y<D5E�w�'2q��?���_ڬ��v{C^^����vB3Z��i�51r [<r�d�[�x����T�9�<��g���@/�� �G��'�D�&3ĘK-��>stMZ>�ޓ