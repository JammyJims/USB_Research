XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	�Z�O���,^���������ڀ����N�
]h��4�)cuSf��J�V�����u�wi�	ms�&q�΢L��t�hG-�i���|��ڇ6D����\q?���P;���gD{�Ț�����k[�%n*�R�C�A�ť����i�K]�Ӻ-s�2����:1}��i�S�AB�`��o2��3���&���Z��'����Ql��[����!��H�*3M��(�ɑI�C��|�Z��v����Ն�_�������]sdG��Q�,|`����?�e����ő�n��Q�p:�"K������G�_~�h1���'��R_K��p@����|����@ɫtAT�L3Dn3J�l�d#]���r!o����W-��3ɒ���|��KӉ=< �B3zQ��9Ũ������N���p����d_��tiÁ�`���J'�3~�hq��碜�lY������������s1	�V��X~3���g�G��_`@sŠp��t�TT?.'�i0�G#{@o�#*��r��3��uL�+�?�1&3,�@b\���� pts�a�ڛ�ף��WfE�C�d��MKAutʮ:���U���I�
�צ��n��7Y[F�>��-�sؔ;�Q���<�7'ͥ��o�%c�)��;*�`��^����l��x�.�ɛ_\y�e�w��WM��z�}/�
�ţJ�k�k0Vfp3S]j�[����Q�u]*����Đ|����q��a'����&�%ǣ17�'�kU���X{1P��XlxVHYEB     e37     6d0NI���'&��8o���B�4�(D�Mj�V�a��8�q�&a-��̎4%`�t��0�酕�rw����h~�l�\`I�>Ӌf\�<�����/�K��c�Di�r'N�e-�#�@@����!�C�=z�Z�gc9����M�OAٙʮ����4}�O�Q3Z������k����JM��?"�꩜��M��C��կ�t��[��Ç�^�z-��`	Dć\p�ԁ F�����ktӬY�Qb|�	4�gf�"b��)���=���a�&m��z�Q`�>���:d��Ga^����Y}�̦�e�!3f[U��X�_�	��)ʾ��-YU|�	i�M����>���v�x,s�Ā�K�T:Į1�kC2h7���h�ABpiZ��؊ήK�M�mY���^:�s����'^g�����6$\Xe,X�� ����[ik�f�t�x�r,E'�3)�s�c�uX|'Ց�� ��`"QZ��CY^h�a�~CO]��|��N詭f�Z4�v��ń!��,
��e���oӸ_Y�D>fu����g��y#��o�F~��E^�\���k+��%�]�I�&�d�:f7���a'ܤ��a�'�^�	M�~+<,
��0�1x
߿�?���K�IGj8�%(=ߒG]z�Nw��4ZA�9�f����.�[*�����+���AM�q&bq����g^E�@���bi�>Ω�+M�� ��M�\��ԇ�hЉ�D3C3걘ҋ���us����vϬZ��|�Ek�&W .���ބo%�����I�+XJ��Ǥ�"}�%�v���NG�������>i�8�Y�g��DBu�ܒ���`��b�cy����G�� U8օ��מj��`�'~��A�(���6En3��+`n�V�߱�� �y��pk'�<��h�����[�����u�I��i�`����b
W�fx���h���Ƣi�0�}&_V�d�i�PS	�� ;��?���`�W���)��L�;��Y��[�2��i�*�L�P1ݔG�WXT�ԭ�l�9#����	t[z�(zL�zS�h�<�;��b�W��V��ƌ H^�K�(6��ٱ`��߯qe�h3�D@a��ė���2G���ˊ�Νjⷌ�5����o�(�~����IJ �1q��{�rY����Է��)<���?Ꭰ��]s��B��Չ�����3V_l�8�3���|#�fQ� f�!��n��ҕT����]��Lw��ĩ{KC�7N�WK�ɪB��=�}�.���Q�e^�[�)~[�B�Ĩ�y���Yl�>Y�̡����G]���^�GXkUj]'��ٲ�#�_&k�EZ��Īh�L�WE���X�U�����D/�Q"
���ٕ�J�.�c�M�֜����,g&��c�(Da�R��AYsll�y�#kNZ�8pw�ą0f=�iq�̗����!�.���BU�[h�^�E�js�e��+�V*%����t� �)(�����7L������N��!Z£�$<�>��YgKg��-�`&sNt���CY�D	��k�zBo�f�|�o����ȃ��Y7L�/���N��k4(���G�%�7$ȕ����9�=���t�]�P�t����M���,�iT�(Bz����"\�����95-�V|�Xtw��� �M.�į�*�[�Լ'��MEOKXb�u�u���5��%π_.ȸ ��e����	����8�O�D}AY�J`ň�|��H�aR�Zeؚ