XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f��8C����Z~�P|!��5.��xƟ�j\;(��	C���14��u�k���:�[�����
K�|ww��Q����lkW��G��$Tv���W"��Q�:!�e��
���K���NT+�5����r�@>���z�h�K���ě�B��.7��g3V�~�ýn�i�����M���V¼��bu��C��㊅Vќ�B�,�Vs�>"�R,��*}�k�Æ���A CU�i캙���*k1e���غ�:�I�`.��Q����:��-?1�)A
����\���in������Gւ��e�f��z��\��R>U�R�_��S��l�6,�q�����Da���'KN�Ą�"��m+�ۧ�h����$ț�[AIkɞŎ\�+=������me{��gH�b͑�g~N���4���f�8��(cN��8�#���.m�M3�:#�_���o���Cr ��a����e}�x�,�	F���l@����L�U���'��4h4BD]/1m�a�� ~�<мpVp!:q�/�=�����ڢ�&V��%(r�5����f_��&*�+ɣ��W]��`���2Է�Kҝ�\W��L�r�Fc��ڤ�&�O}�����'�2��{p{�Z�P_���n@":JwB�K���2��/������j���l
3��S�;��#���⭻���1�h��}��ƌ�)<�z*���0y9��2Ws�i���==��;+m[�%��`RRA��~[<?!mU�TԂ�;	:��vC�zXlxVHYEB    6015     ec0�n$�y���zV}NF{�R�=�9m�Ș7Y��]h�>s���P�G����B�n����X�KOÕ��G�1�0��1��6��s�y?�ӫr/`T
X�	��4?��`�:���F0�Z�F�;tp��j7�@$�)����i|y�������S�E�`�/�XG���2t�_1Km����� e�_;�j�Hds�(. ��P��=��ؙí�.ݻD�͇l�J4��Ոz����*i��N��uZEr�O�j�Y�9����ա�
{K� ˉ���2O�G6Jl8��b&�w����`āu�srt��Z��-RC� q��������7Z���"���9?W�w�U�>#�d��&dq�v�\W�傾��F�8
���D�/Ӱ����HC_F����9�
cI�,��.�z�.��θ�s3�!j�í��0D�iz����}|c_�BL�9��i�P�s/��~�5�>��l�Ḳ�:�_{(���>��l'{L�[��}6�I��Cӽ��&I�� �>��L�G�j��jpҞ���z��@0�9���Y��X���٬늄�&��h�F�v�τ,������ �o@\����Z�ʟ3e��r|��Ni	=�����s5e�������kFǇ��$����(@���&�?�&�ڇN2G á���-�~}�JGj����Q�H��dr��Fr�� K�Q7$F$@������%�L&><�]��n:T�����q1�0jYX��O4x/����S(�x�y�U�P+���4Nlo�v|�(ɨf�PP�YF�i��.�)� -SA�v%�jȎ�A������޽Au�T�����nc�а\*���SC�,�h��8�|)IK�&L�������Ea0j�#��Q jL�T�XǊ�o��!�=O@�@MD߈���jt��J�Gn��yQ�Lf�İ�r�m!<)�΍�$�ʄ�y^klHa0���kKώ���<�I��z*a���8���%�r�+l�`ic�Ɉt�W�S=���G@*�W��3&se����S�5�EU)ޥMB�~�,�e��q$S���V�P�˪a�E�(�랊�|RFX�\���n���9�D���&��n�h���RƲ��
�,�E�:����{l��E��Cn( ^��1�.��D_m��h�Z�һ'�ȵ���x��Ds)ۛ�ZB����9I��ķ���t�z��.�u����QP����.Te��pIC�?��6~/4�W G0tp���l�{R'��{c��K��!,���/~M�#�?�.6��S�2�lF
DB=wy��p�/A��Ԝ➗N
.������]����Ğv�n`�.�N��wm�vr��[;@�rS��	F���Ff��P����~�i��=Ֆ������Wg����2�j_ʅ$*��Y���i^�Ie.�R��.���q)7�i�����(߹�2%��hF�A���O��XԔg�Z��1�{_Ղn7����x���wm�G�t�~���ş���@�1=�c�W���Q��`@�b�_O�)�C�/����o�o�[&6��Vl��Ʊ}=�uf��*�}u�`��{�^�P��Z"a;yoP$��=�p7H�{ntH�>4y?g�j��jT������Z��wη�!㎡�-�>��:��"�x2{]�7�A��f;i��+1��3��k����3�̻T��k�`�����_�$i�b  ?�\M1F���K�bU��Z�>F���OĪ�
�k#���c۷/�	�n�U��d�����"����S'J }�t��`;���U*�e�ȣ�o���F$��-u���T�UX67P�~B�)�AO^mj�N8�Y��P��sF�� '_"/�0�P�v�h��1̏!�P��/���+�=ݳ��{��.� f��y@����!K� 8jH�X��O�޸F��F��I�3���Mhh�<Ϣ���&��j�ҝPjB��bb)��\����� y�|���F�˔��f �M#tζ5i��ϐj�0�B�E4Z)Ğ��s$�&r��𢞜ޞ�Y�����K���-R,$�,��<�<��u#ک����=�����}��$�e�
��{�ȸ3���n��I�F����w���4�D}L쫘��j�/�~J�p[Ɲ�8�����3mV�B�a�A��l�h���$3WM�mhGc���Xf���?ǋ�|<L�G���K\7f;`�~��)K����6X�|6P��$��}��	�E��)ն�)�5v��&���}��b&�����8��#][
{��|�#��{�i�HVBɒc����.�@+���
t����$_ ���-$v@�æ
m�A�28�U	Ϳ#ŢQ*�� ɳG1ƞ��x�c���
N�������,bk���#T�XP*�"��Muc�T��K��%��$:�q��	�t�s&� �M"59=�Ke�پ+��ꊜ��&,m�^��_�i��2��ݴ�9j�w��G�셢��:�я�6�k��74!P�C˒T{G�Dz/�ЭSb��6ĝ��_��ZK+0�<�I�L4�V9�8r��a�Ś�X�z�+��+�l<W�5�C޻5`ڤ�.�-�O�]��C�hX����R�-��#�q����?��T]���1;����b�?j�?��Ŭ���_��������M�6�d<f�s��2��FOӻ�8\�[HL�(��o���Ζ&e�ac�&�A��i��?���ƣ�G�a�(3������Ӻ��WΒ�kVzI�M�Pp;C O�=�9���*�
���D�M/�{r��p�d>��n�ZÂj�����jg�k�[&�V<H��O���٪h��������I�r�=��F:�?.Y%A%2WEС�d^���{�6��eؐb�`�L���	����N,n6��Y����b�v�G�������<]?3�]���WdJ��7׶n�Az�7��+輺u�+�kڠX�H
:�%��a����s���:�3���r,{�?��Xa<����e/�8�RJ��Tx�.��$ԅ⌿����Lÿ�tQ1OuXO�n��%@!��T�l��N��?G���(����"�}(o�"� � �b��@�E�r�$�(�'4� IR���ӕa�����䎸�l6NT���zo�� �Z��@�9��.�ً�!N�����K�4��f� R9R�s_�VAG3��UN�nsv�T���%�0}�m�/����4�C�[�}��h�^�xC�ő��/�!`1ht!
R�I踥-,=(��"���BY��d�9T=K_0)L(�*o�7��Liy�ֲځaTk@����`QitQ���dU�kz�؃&Yţ��=p������ɞL��l�=;s�dt�ơ��X�R�s��W� �����a����S�t}J$���r����J��*�ع'���!b�o	w<fR��l�.2�T�^c<H����BH{��G`�Z'u-"W:�9B�au|q�jc��ߺS�M$�#�F���^�C�ƽf$�6]�.n�PV4�yT>g$���h�f�⇾�4�e:�6�����r]	v��J i�=t��M�祙v�Y�8~z�#���;V�O�yZ�qNvBU�9�H	�$,����9a�`������3����yVQ�@�'j=p�d�E9�IO�^le��n\*���"�����VU2x��C�_"������R��	J���}� �E���5�j��