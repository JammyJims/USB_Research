XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7'A2o� _���u����7��V�h���l*�p��d�eP�A�T0&��G��U�tW�`��Z
o�=Mxg�:� J��"_^�CzM�?�O ����q� K������>7��X�����us*8\�ǆ�Lb>�bB�?ׇ�`��WHɖ�h��Q�>N����r�_O�u�Sem/}!2D��1�N7�/̾r�萸;zcȀa�]`L��픘{F-v�:
�������hNm#�[���a<�S�H�5��%i�(JBFB�Q�3u^��gG�`ٮX�:�,׎�H����~@�:��\֎�/�����S���(���Vc�c.v$�~����p��G
�*,�
Q�RAz-5o#�O��nϘ�l0Z\�prz�th3B �%x�u�)�g���[� 5�^�^U�D&�v�t��F�e��hU��5Y��>JI�L/y�i�a$�ʿ(ZǶ����~K�"�H�Ph
�x�0��+IcY��L���Oɭk�"���V@O�	��9������}�|c����R��<���8xs a�Iy�I�s�[���T�t0��leϽ��kd��20��&TI&��W�sU`ǶԬ��·/��B=�XȲ��e�����h�߼;���G}��Es�^t]v�
kA��(�Zf#ZΟ`�%<�^j1~>��=�V���� ֽ��)�G���������Ը�e�~���s�f�̳
@œ�W���[j�핹��LP���g��w'�����;�'{f0͠;P�cXlxVHYEB    768a    1930E]�.!�����kT+��{-�h��q�̑%7<��͸屲�e��q�&�O7��HZ���P��(2�P�V^v���埞�kk�h̹�7��!��Iچ)l��"�y����X�������;�|e�]F���~�94]� ��pP2Oh��BtK�as�嶃�O[����	�1x�>C[�UH�E�Ga?f���F��2�)����
�iE]��p��R�W,�J����x��OW�*i~ﱢ�d�ك�5Us���(�*� �>��������[�~���(_�������#hy�[���^�8hi1�#�O�bN�T���9I�qJY%)��mM9�3��ǩGj��??x�:F^ޟ�D���(���P, V�&�)Ƥ ��|!�zQ]���l�UGj&�N_��9[o6���{����:V�
Vp8,նEMV�W�J����]m^�v�)��a>�E�m����;z�OV�����	l�C'�_Glg��kK\������_�t{ڼDO����g�u�g1���*rwI/g����K������"��i��:��\U�#;��f�^?�R��qfI�{�{*��^�a������bh/�G�Qe�Ǟ�!�zR+skr�n��ףv*N|��2S��o�=S���)[z��[���K����e�w��~tE�@��2�@w	�e޻< J�K#��V&�B
Ԣh(έ�Q��� Q��D~7��\O���W���
$$��x�S�zvi�iN��+�]��1�qZ���V���a�yac7t}N��4�VWX�T�h�V�vS�EN���?M�¼�<�:&�X���$�"��u�A�^�K�����쥂- ��q���/[b��ON4�X�����*������e3�Ӛ��|��W��[q�[Y�,�[|*qX^�d6�ػ�D�/T����;�B(s���W�|��*k]8�:?���`�YM򺓓bm�T�R�D��rD�苗_3dVQ�P[�;���㫾���4u�"�d?+֓�M��-����v�D�0�&�������R�}V���l�I�i���4[�H�C���]���$��'zF�҆�w_8w��<�Τ:�g�y ��;�c7�F=���{o�v���!���@�fe��j�WFK+�hM���ho�ДP�l ���o��]��#�S����im<����P�V8����;�S'U��\����!��l�:NZI�����lV爤uAӊ$_�A����Oԟ;��0��C��l�R3�����cW�u�9x,/,A���M5����U_�g�H��\���0A�Q�e��!��v��A�q7�9v�T�W�ꍁ�F/߁��È�1΅m��^��}L��KyI���i�з�i���uRu���)�K�S��х6��W�%��_�䢯L�O����'w(!�x�Ԫ��:�s �w��8��"m���QoH�@\���^lib{�2�m �4����U�Nq+�ApFc�Q�S�T���g?�)=�0R�H4������w�A̪s�|�:I|���Z�n�d��g���yh��T/F���H攵��B������8��딹d� o�ֹn�����f��'&.�E����^ ����0���Z|=~$5��9ܿ8��0ˉ�4���Q$�Mj������]�z�!�j���HL��S�h#�����)1���\�g�L�&�.[|��u4���n-�������F�%d%�w�N�@]�J����, !ZB�Ua���P6��Tz1���B��zh��f��iH��HC6�ǳ����7n�XY��$���=S&z��)bu�/��c���4	�2_kw�
��5�(���%Jx��]���V%'��WS8��-���V��r�gșvȁ�9�����?w��8)�Θ�%0�����!�� ���:L��F��4������x �$q�;�-��y��ٹmuD��d��:u�c��������).�TJ�`hmP�QP�N��obl`���w��t��P�~���-wM�l�����uz^
]�/t1��z��IoGR����#�[�S*��������3��pJ�?���V��;Ԯjʽf���Mյ����T�C�sA��uB_W&��8�9�i����5��αΌ�C	��{�&1pD�����Ҍ�K�%,��'�߻��k��.Ǝ��k��#���b�+��[ZrW!�_�@An�zw�w�K�>�E�(X�/3�/����S�$b��oΟ�5�X�5�|׃�w�TiE��Mli.%��!��w�[+<P��.ڠ�B$ ���tow�a��# �*�i�s���]A.a�v6�,�&�u{ְ���O����@}��zu9� w�C�q�W9�i�JYV^��ʮ���U �?rI�n$�X�vb��fR~W*q���ƺkZ�b���m��޴\p<a����zS��V�^���Al,�\��ﶀ��{K$*�`>}��� �FkVs�=��. o0'��jb�u%��ۇ?�w\�Ҫ��X-�^�Ay�W����ܟ��B�\k����輟�1�Y7;b�V���W��H�L�:�@Hsd<�r�<���1�R�xu�c�����[ ���{����'<�c9"B��w)�ë�J-~��FU��!��b�R��g�6���5���<� Ȗ���[�V(���z�C���9宊Qs�}���w��\��H5��Zfc"��ŋ	]2C8a�\�|�>{������竾�q���/�S���;KW�����q<�&B�Ns��(1�6a۟��#+���$A��l7dao��i�*iD9aX�$�U�˩���7�5G��q���t�D�0�iz�+2Ϝ6L	OX������b˃1q-/zy*�w��$d�r�)��(Ȑ��fJb�v�w�<�"���t������Í��8Wz�W=/��	�w�[
E��K>�<�3<�H�R\�0��gfժ١�;+�zו�����}R���R��\p��R;)��<�,Wp��X�0��*��x���O+f�Թ�0s<��<
fC���#�$\7<q�h� ��Ch��ҧ�V��I0 s�Qyk�8W�8�� ������4���Er3V̾��0Л�T˥��1���l�����$ ��<�	#a���"XS(���hw��/b\�
�,\���[6Qcf}>�`S�{L��{`���;ڏ����a�*>���®"�0���3ۆ�Lc�q+kΚ�1H	ebKZX��m�zdK�I�
��i���a�wB�D\~�%�y�Li}-��z���W����Q�L����h���<E-���InL�\yM��3�B���B/��~m�f�BtP����)m�)5�\�nuL�m�?Ɓ;Pu��H˙O��_3ł�J?��8���M���Y��쳳'!���x�P�����~�e���-��MK��ԢJ@����P�q���o���
$��J��N�{g�LM���ׅ���m�Q���M��St�J���$e�����yHRu�
�IU���4'U���f���&���[�B�~L����C~X�sr��$�9ccV��=6��f�����:����vI�+XM���XLq��Z�?���<6��K�6�%�9��eQ�-0y�ʓ��oz���Ls�e��K�l�\,n+gO��M��dG�k[Y��(O�!X�ɸ>�U���ț)*b�!j�A-	����;܅�RL8�FD���<��`m#��3��Ύ�;���������/<��X���#�)%\����5����'�:��^~��Kn|�9Y!��s_�5�=���9l���L�ӊ�ť5g�f|]=e`�ԡ�\.���~�R��ⲮB�����t���j:d��=��L@L6�nh�0�=�q��<z���%��a�h\تz�D]I�4j���h�v����5G��b-���#cj����b�	�[0_���͇&�l{�.U���Bi�#s�<�YhL� �m/�;��x_cB�3��<�'��H���hFݺ���莓k��	3d���n!*�
�@�~�5��
���OR��jK�/V��r+���K�-���u+�4��i�K����~�M��ՈO��w[4��^��LӦ��>�>�#�@�u+5���Yu��o[�����L�o
�ӑ�廠�
P<��S��6�mz��I������?��������JPA�}�e�c[��X`�&\$&D�L T�Zh/Μ�J�u���혙�+�3۽Pp��nc]���O�Ge� �0�	��M`�ln�W�_�0�G���q�N.����EBޕJ��N���[�Ka{4]�sFED�|9hOX��0���r�֥#��a"�P?6	��zA�� �����%G�s�����s�1pN9)�o�ju��}Ѐ��^�šw�>�_~���`�^èZug�.:C�5��yA�8c0�u�˶��;��X9�R*	l�J�ۄ8k@�����dL%�����GCW?Ϭ���Sւvo�z"����{�,x9�_�ޕ�ˢ����Q��h��ވ�fpw�S��T7r�����/]�����.����6�$&W��Z�}���������D�-��d����'�d���$�L�bժ�Q>���A��$r�k�1�V�pمow�k2�߾�x���W�w��O��D\�kX�=�7�T$cسL�����ل݈�-G5��uNZ�c��
&%F��R.͋��^�=��o~e��aakC�ޅ��$�`�'�͘\��eˋ�؁ئ�-y-\�z�>�"�4��)�R�G��y�>�-�Ye�H�O~X�ȟ���ບ��O3��PJ&s(W	^�64�n%���6�;N�<�B��u��a��t����92�'%��шrf����#���@q��֒�����Ÿ��g�A��9X�-��f!�x�s.ýR�Y���a�&��;uj���pR��"�3x�2̤M�E�|)�/�V^D����2p��Zv!�����ׇd�������P�-oJ������[6��ejE��L�&pni����E9fC��g��^y�g�'���XRW.*x�E�:��x#�b���N��꠼P���7�cؑZp1d�8�_�v� iAW��8Ƶ�ζc�s��!��t=��K��3��V��ӎEJ�$�U�=�!^�9d ��Q�"c��ߌ@�@�$	u�D���"r����t@{SpnB5��\?������Jt�TuF�ʂ��
������Z��`�R��"�j�L&�\�I�U4�"%hk�{jzx��I �������",4	\�0���5p3�6ftgo�=v�#���G v%T:�R��7 ���adɅ0�wU�����P7�FéG�����3�v��2�ycd���
K�a��{�N����kM8�%؋q��r��IFX~�Z�[��?$,w��==�Q��ͯ�>C��=r���{���������{4!�r!p�j�3c�����U4�i�,,��eD�����1X�E�o崹 H���B_�Y*�)M�C���v�|�R{CC3��>M6u>OH�m��Y�!Q����ݪН	�i;&-�a��?Ş��V	�XO��Ɛ�N�H��ޣ������^�G�A1�7"s$��l�fH�z�=}��J?2�0	a�l��,�(5 �ɺg�1EC�A��z9^8m��=L/HO+��v�|t�Z�kf��ɔg�|�v��(�7�<�V�S�����`��Q����9`��#�|�ex<�`��^�Y�碑��E���Ag{ED��7�g�B��\Fj�/N�с��pt�R�V0je���a�bfW)㎮�}}!�Ս
��� ���	���V��p"R-�%ئHh3ǚ�g�#�����~�5;p������7�̈qN~��-��	�9A�i`?�5��%�9�-��{���"�ֹ�u�WD�ƫ4� N�3��`\ȁ&8o�>��|�����A������_���˕�Mv3q�߹0+��)x�:2����y�/�Y��:�Z����΋2L��N<��ƽB��Q��_Xg?���:��o�a���q�9����A���`�����K]��7�(%������?�Q���%��¶662�e,��s@-V���oyB=�B#���N�j�c!4�4�`ꘋu#D���2C̠9
`)������~J����Z�7F/)O�'�f5�k���c�/>_0F��S��F������(5c��D;��cH�H��P���ִ�?�'������� ]sW
���!�� l;@����w��޺�!S�L�j�� #Xu�Ky=3����rfc�����m�P>�#l7=�	8BMfݎEI��4