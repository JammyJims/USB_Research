XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ih�I�=�Pq��b�x�4`��i�4�_�rЦV�ġp�P��Bp��o'pW�?��kϞS��mVg�N������V��ڤU��M�>eC�'M�|u�:�aAy�� ��]��5�ע�_��O�-Tf�&'���G
it�g���Za$�:��<���#'Ե��gO,l<���ŏ�?��p�J�E�)�s� I�������c��C���X��n�����O���Z��%��AC� E�>�E��Eq<����P�=i�w�9y�C�&���/��21Z�:0a�V��$\j���MЁW�@�H�}�\�>¥VdCnd4;�m��ﾴ�XN�V��a�քG8.��W����9��f����������Ɯ��;6`��^*����P��
>̚��E�LZ��%Ynқ��4o#�����#�z�:(wj��dQ�t��)�u�l�#�T`y�DHb}�Fo1�0w�l�t	��=�W_�gPŐ��#��m��*�G��X�`q�;�I\�ȴ%%\ql[,�+�IC��X�t��9�۵&����S���oߑ�u�M]�L����B;-���hbO��3�A"w����(\yK@���"&���9����1LW��趖A+���,]�w���W�=�`��=O�0��u�I��3��m�f�\s*W�"���OT��h9�߽�����5�� �G.c��X���?����sA�&]
���}
0�nz�A IR�愥""l�d�M�R�	��hC�x/���XlxVHYEB    20ac     b60# � Lr�p��{�Ⓦ��4@]i��µ8�3����T�7/��
�j���s<�/�-3��s��o�[�곅�iE�3q�6����ڤ�N~k^]L����|�MB���X����)��SB����> �>03 �ZD�q��Ɍ%k�R�3��J+5�X��a����-�n�G!�H����j�i�.S�Q��m�p��%���&�*1�������7��ϵ�zaF�{����}Vv3�>�����^�j ���T��_���4D�&@�[D)o�&��S-x8s��,�Ħ<��׎�E���A��zϝ���y&%�i5�ܡ���H�e߱ᰒ'_;Px��٧�?(����,��Q��Ur4�\^`Ӷ%~�Q��ȶLoy+�K��0Ƈ?�L/�s'�l�;`����3����O����hrI��A���6�� ��ނ��M&�`YE"}�y�Uf�ͣ@�U��ԅQ�BQ��E���l�u �Fj?"ӂ~�K�)c���J����^C��F���0��3�	���z!���jJ8],���pN��������T}�+a�>o�"�s��<������5�/��a�!�t�Q#�8*N����-�L�6t�ff0����ƱC��jRR��R<��0���D3���f�>k��������U=Z��WX7gW+��_I㯆Q�Y��e���>O���� )w�sya	�o%��>B���X��˥�mv�XCr�ߙQ��ptV�٠�Ut�����L��IZe�o��X?��ݷ�K����	���n�v��X�-.踜O��Ic� :�#��R�'�������������-[�,_'�9da԰�m�1�����ɇ�ff�T@�r���rC��&��@����i�� ��Uf���(l��P���*x��s��ƀ�P1p�J"�#��8��9��{��<T�+\�٘��H<<�y��V�k~}�(���K\L�͞8��V� ��;����̟���p
�I��'�E�y]�9/03��:���vj0
(��[���a+��s����Wt�S���j�W�`��7�}6�a����#Y$8�Lz�u�ϽHY��ya�_3�߂C�Z
��PT�5�� d��̏��咘4��^����Ra��Q `G�UCi��My&)9�
O�r�]JU<�<��ؙd�̽[��w6��~rE�y��Vc�M\�9X��!,�Vg��2�u�G߀�=P�7�F_$�xK�:��F���
z	��yeY�x*�!}�2�M���ꉩ#�^.�$�/����}ٿj�|s�7��=��&^J��kn���F<��@�Įn���%�5��ug�����t��ˬ���_�2B!@��ur�,��U8*
���H`ͦ�'�Dڬ��~��<����Z�7��������+���A+�du-�t�2�SX`s���"�8��c�ZKa����JP�N���`�N҆�Φ�U�W�^���E�N�,�D���|k��K���gp�A�ǣ��I#����g�	F炁�����=W�x�H �gqp���6�Q�/ӡq������v��R%���[�s�Pf���`*��d)4c/s���(�����O�����`��j�zoJ�8��|��p[~�z��ݝ�@(>���"�\��u��¡�����G[b����J�)���L�n�g"����č��f����F]�Rme��MCF���$�U��B��I�l�;�~�⮬��P�&�����F��m�7�TdC���D[G)<w{�=�Q�4�yɀ���]Z��O�O*��`,��pZ6�<���Z�zYz;=�����N�H��LcԘ��/K1�m����%&y�L�r+�N;�{�[�&p���-�ߕi�2�����wp"�v�	?��i��F��z�[f:��*��ҋ�A�H�%W�dy4�2Fr�/�4�7$��\�	S��:w*�B/��ˋ�;ɸH�~���E�kI�B�`~u��y@�t�b�ݸʏ���6oJ�8t�y]�(�ɷW-��(�\��g>jo�H�aXpUMŴp�#��P�k�}	-�/��d�"A)q���5ZQMT)�����m#@�d�嗉�0 ���vU��1�'�B�/3�&@&���Uv73q���rR�F����v�6T�G<���<���F1�!��L�P�(;�4��EZ���FMBL �9"�f��#����}�_�Jq%Y�Ӈq-��G�Xk��;�i�]��<�t�b1+}IR�N<�Z�m��x��wX	�
+�IS�dHA=:�` EW~F���g�eC�yp�����n�y:>�3��kt��n��

�>v�YKL���b�����u_uCy�2/�6���:���n��wv]�;M(�����=�N��c���``�;Ʀ���BV���vwn�f����c0I�XU������N��?�	H}[E,
	5�Z�eQ ��'������z��<�f��@��	��f�Cu����J\}�P6b��H��q*��co^��q��ȋ�`M��-�ÃgS=��hD�Ζó��Rq�|q|6�>E�P�s!��i"�
y��f>���x���|�p�]���O���p8:��֚���>�s��;*��^�a����3Գ6Of	���7U{p�M(����\^�F=������<]����Ɏ�}^T���#�p���B֬JW�s�����.w���9�b�X�0T`ၟ*$p��ʖ�q]��V~0�
a�V�J8cO O�*�	�^��^�@�����ex5�"!��'b�$ã�NඩU(lV�#a�3Y�)CP��.�>���*1H%�Q��F����ţ=�s$�z�>�%DY⃿io2m꜂A��M��q��;�r�!U:����5s�!?���:����"