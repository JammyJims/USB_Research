XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s��*��c�C����o���!7�Ik�R���	�ӁL��]ķ��Λ�bQ�k��g�Jc��ƌH(��0{#}�����t����8Kv,8���|J��r���h+g/�����r"����c�US�����!����Vp�L��j}�	�l�M��+x�J��͠��E[҉�R��v��G2P�q�㿇�ѧZ�v�����Vd�2y����� �Q*k/5C���jv��K��Ig��m����0(���m}�/����n!��ͅ�سj}Z���ѣg�<y��N�aޮ��7����Y����!�Rmڈt
�t]6��k�r|z�r�k��PZ�ܑ^6�^|�=��_Q�H��������e����ZJ��A��/�&�N��Ơ1��G���"Hvy���Z��>]3���X3�4p��S$��܅��(
{>?�nO���!�H�2Q )��@g����^d�Rz��Q���J��o���I�q����VVd��ig	�����D�_Ӊ��Ɩz�����n���>�Oz}�g=������&8���z=>�e�n+�f���7����"Z�2d���wۤ��e�8��SX֣����[Ҡ/�M�	Y�] y�pj�]��)N�2������r[���5��m���Jg�p�������_*���~e���a�����[l���7�Ə���$t�a�+�Q��]�3�'_`����L1r$��RpI�� .N#�&��ތu�[_z�f��~ٿßT�
{�E�v�����XlxVHYEB    a282    15d0B�h������}m�lf�����1�����Na�O9��ɺ�[H����c"�
qM�1��^9�<y����s��5R�]��u�НXfu�Ҳ��$����q g�D_�<&7ȫ�Z
K�.�Ėv�b0�/z亐W��21vsKz�� ӏʜ�YV��B<ܺ�-��O,|B��Ɓ���1��8�$P�$� ���E�5BR���Iu=A�5_?p��E&BN�ǋ�f�uA
��--U{/eSL�6{9�.��v
�2G������d\��d_�Q8���`R�b�h->��p�<�]'SVr��5�-�\�(�ɇ���`��?+�!������a��w�*�K��4��5Ũ�� Ӣ�9H���,%3��&�ѣ�Pd��!I��Nڛ��G����Y$%��6�8�Բ�5v��
�j�"���)���Lm�V���uqo��ʛf����gL�K��F+[�*�끷5	��S�����ĉg�*�6植W�&�= fu�5���b���`�~F��I�BBwe��U�s7��]n�<��9'��P#5�76Yt�j��)�0{R|4���'�Y	VPj�V|S���B�
��\��c��^G�g���֕4��?�3�jI]�|��\��-���v�7{�oA�&�L����L�_ N�2�w>?�c�C�H�>��x�f
�G1 ��Ӡ����>�S.�V���z=/�Nk�P�C�m�C��'c)wFi�*���~��$�2���8�##���×.��C�/�8�#�M������e$Ӄ��q�ihW(Q"nl"d/W�86a}"�T>Py�]y�<�/�2z�p����%�ٛR@�<'+�s��)�Xb+f�߬#�r�ꑙ7f�)��EՂ�iy�XP���;���}zq�ܖ��d�?��ؠ�Ckl��9S� �Cح�pI�)ix`�b�����e鿢��o��ys�P�h�"�8�kEPY$z�ՙX�I{�#��6e�7X�@��ֽ�oIMם_oz��Ҍ�4����x�
>��"���3
rhR6_Қ�r���H]e1Y�,K����۷�(ۨ��t��t�b���w�WS����N)�Ѵ�^a����M�yY��L���x�FO��V��JEO�<��} 6^$����Y{x(#�D.9�=�?Ne�����'�M�����s�.������>S)1�[������7�����&~��)H�"s�3��P�'2���Y��#{�
ǲ�Cg�K:�H���K�FN�x\f�6�[v '@�����څ١c�(<o`oW":_��8�"�*��Ŭ�z�Yf}k��1�������!�`P�	I�S^��t[�KZ��S�:#��ƾ�[�D�""�w�gb���].�d�k��]���En=7L�!�����vf��5�u�႐R�d"�q�f���P
�� �X�H��TRI�30��v�XZA/������"����L�M�hl([� Q!�:c��|�
���d�9��S��WK�aW�
���BUn�Tݬ��H�R#���'t��
Zec�;y�3�1K�?�Y�G�5i����ī䔔B�Z��S�#J�v�hp+K��s�zp��� �&���"T]8�$��}Ȁa��y�����zvAeJw���?zk����;wZt�I�έ��~����l��ё4��N	;���Xa�DU�#Z��K�;�ǈ��������{�6��g�5I'�
0��@����H�,����XC��VV\؄��8D�m'?	�ۯ5T�*<��zg7���5��mu��9��l�"O��
�D s�/��b���<x�D#��޻lf����6{![��Ƈ��	�f�+a�%v��6�-cx�Sݨ�kϊny�s�����/�GƇ��8�X$��.Y�{vX�(km\��,nP�����D�ƫCAk���xo m�J��7�m��x��9 �oU��#M�@D8�~��ɾjs��^�2���}嗪^i�N�����K�\�^��H��E�D��-$��R�2���R��!�1���M&�]��qP�M�1����ч��s�6a��À������`b�σA`m�>F��N��G�f%+�wX�_4x ��gʺ4�rh�̇^U@������5��G��R�Mmt�F-��*5�5ڮH�t)�ݰoQ�ϡG��5~�9�;�-K���(Ez�v~B�_���V��C�*��v�B��~Q��Y���L�ЧC�`j^X6зiY�f���	��*o�+�j�QA�2=h�9��J�[����]/���L2ϕ��c�%_�jG�#�����t�5:D,����h�NZ8�G^+n���T�K��ߨ�Y����O�_<�GDs���S�<\z���9�p�� e����l����E����}.�F�p�~�S]Փ��i
@��SҙEo���qOy"�l�=68����b���(c��%K�ƀ}Q�!8؁WM:��z����B\�b����s��~]{�+�,��Gں:s:�j��'"�8�����^���|乬!��>�|�h^Z���Z�r]���+��z���(u׾����e�Xl��D�9���~^�n��r�L��%�叁k*���
*�r@�Q�6�uҔ���!�l~�d,�e�Y���q���9����p	�(� ����w�����Or��|������W�N>&��y�����:�x��t�e}��"��ҒbI��\�ew�e*^wt�P3侮y�^���B�/���j���=-r��·nG�XE�&�H�]��P���E��m&I��Яڥw�����:�W���5�/H[cTqaj<��Z=��L�^�hl���_�Nmx_U��T���A�q��]G�����Foa�)g�,���v57>Xfɥ�(��I+�F�xJE���9M���۠�]��*R6�����\��]�Vȩ:�i��:E�����ゖ��rf�J�ffĴ����NY{r6��	�ݡKs���}'r��¡���~�a���%E�o��o���>�(����Z��^5��'�9�}eЄ�~|l��f"�EH��\��\��;���;����e4�s`��z��v[Z0�;.o������&a7��E�dWZ��Tѹw�&0/d��]=����F��UM1'���6�O��	�q�돨�1]t����{�i�VLR�k�hM��h�93@ʼC�Hh��@N��E1}�|����Q_����}���yFI�l�S�!\N�G��B]��I�:e��`+��8�v!���Τnm����/� P��}Z!vOR6x��'ϟ��3KR3a�8{�ц-�b��()��z?ڡ��,�{נ	[��fݦ���1�煙����Xn
�JJ�q�4fZ����7�p�����"�*��d�p5��܉}����t]�O!�.j��Х��C����q{�wN8`�EX�Q���Ҹ���襤g��]ⱱhO�&�$��8�g���x*�t���4
��y^��l�*��yԅ�M�32�&���9U�J��J ����\�@@�o�=e���ո��2%`�t��Z��ъSnx	Hݼѣ8�e"����ɃEj� �������pd�6���A�v�L+u�+�9*�Z��|�G�4��rǠ`.��p.����w|b�{��N���5t��Y$��<H�De9JBq�E�򹽳�.�N����N>��e�'����t\Y��^�(Q!���0��̐�$��O4��G�<�|�{��S�&���������}�t^V{��P�#M[gl]�P� 3��b��s�]��mP�Y�A���A���s�"tU!�c�{K{b��YD�[$�ۅ�C�n>;��,@F��\1�%���$N�\����r�$�G��������찭�>M�BK8�+�(Y9�4����!�G���Ww����s�F�ގè��\K9�"3r0��2m���.~�.-ē%�@F�J����.HL�#����G<�+����,�$V?��|�OMe-W�dЏ�Y�S"��@Z��Иjcr'8����q{�S�ߔ��Aw%�ӧ!���E�T8Y~�y�O�3�m�x�u��ώL�2���@�4�ך{)��@."�0:<�e�"��������U�΢�&�ڏY����a��r�등��p�io����<��������8�4Gt��T��������a�܍����]��#����)���̿S'��+N5�	땙���s���v@�
���'f|]aP���z��ö<��~�wv�E�w#-�P|�@��?�gg"$O<��Y�p�}E^��IA����;!FА-�EMj�y���4�x�ڼ�r��}�.��S=�/�v��hr�C��-nh[�Aq�Y7uJ�M�m� G���ѩ�H�􅆮��a���7U�LbL��Wd�z����F�JPQ3� Mo���}���������Ԩ�O�"��<w�^/J�`�����[�|�/�KQ^�9�X,���r��W�[�)7~�6\Y����ƨ��n��	D%�Qw���zT��X"j�y��nm�A��et��N�̅�g)���%��L-�
��A��e�� ����F�[A��X�ζ2��q��<xO/K����yWM�(o5��٥��*d��d���4��h���+Vԟ2"q�����mr�9NZ�/�T�q��ȟ���6��?�4���Y*W���\�1���F8�>j\�U~l�x
k��%�6��Ipak�2���[7�>=%9r1+�:Rwȥe<��Gs�ķ�a��G��ӜF\���3����ak#愖���
�U<����ey��dq�[�����%Z�[V��)y�^(��ܭX}B��v-� �RY/Vh\r�?U����M��?�)+ubg*l�
�+��)���8Q�R�K��Ԧ�l����Q^��0<������̩A�&���iZ��x���r��W~1�d�\kU�ʒ,ߞ겭��&�h�_���7�Q�.��| ���VG���
�&o����Edm�j2�;Ƣ���0�oY[��~�v���i5a���|�IvI0l�F�]�p�����wr�����������QsgZ&`��|-ir���*]zl	���ҿ��|�
�R���f;��$Q�v��^��߫����'~����m����8(�iҨ9���G�d,�p1d�WO�Uʙ��A�X���Hܟ����C�HH��V�4u��WA��'`��A�|�FQ��+H ɭ�g��Os�i�x�]�`5w1�W�*�TLF��.ui,T��QL�B��3�u�N|��Eƣ���5�ko'�&gZn�Go��oS��RU�y��f!r�ח@纨�d���^�V�9�Ɩۛ��0���-���N_gm�����h��s����Iz�*�f<���*#]�;�>5/W��Ь��]�>лv�p�lJ3)#�9E*��'Vp���c�h�j�ߚl9v6c~���{,-^Q#bڍ���β�!�н޳�S��J ������b