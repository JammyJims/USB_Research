XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y��u�2pVd�J+{?�A����*���ͬ}���(�z� ��p��z`^���'A����M�0{���F���%����7	ƃ}��_�:�y��8�E��+���G��>�3d�Y�M�Rz�A96�����LIP\�^����7��irs���V�и�#�mR0�o�o��)�R��O�5�1D��@�O�Y�v�D�"�/z�sG��R��y(w6��\�`��X��r��I�H/��S�a��|#/x'���A}��x��8�J3�6J�d��O�1�}�]����b_ x,�>��E����Y���]�b����i��yw����w^�4�5ͦ����4���?:?(Ї��:��*\�)&�q���e�j^�V[r������̒Å��^� �ꉯӔA/y޲P�����EM�����T�K}J����_��ǩ��r���_C m���Y/� dLV)���eXƮ}��~�4�ﱋp���.�PC�$���'��}�����!՛B�͓V+g>N������ h�)~�\*����x1(gx�2��=�pd՘�#,6��'��Mܼ���'��!���� ���^"
�Aj�]*!M ��Y�4�@��H��LOA�����w>�Q���s�OB��S7dNSE�$z�Fڹ�[�SE�00��{��vb숖(�o�w�e׃\P����Ye�S�R�����J*e+O�M#����+��4��r����/�Z�"�ͥXlxVHYEB    3ab7    1040Up��u��Ybi:�T�S�{_��s����ͳ$'����#<�ª�S�;�M�=R�\�*��7�����f~D����8%
�Y�<Χ=��=��l�o�Ӟ��X>��Ư���l�h��T!M H�2�I�d�����L�� ���]�7��<!�
Fփ�?J�A�R�=�VP�+�|�v��_�-"���@�݆]ϖ>�&�)i�p[�}������z_z��3k��:�. �+�v_|Z`:^�\ch3��;0&Z��L����u��[Z���E[�]���3��D���b-SEn^���7t�1xp�G;�}�+߳�����m��c��
�:NpQ~�R+	���f�\P�>	~�/Kq�OE�ʬa!��`Sڱ�~t��B�3��(Ԫ�?��Q��z��S�)�Y"z��8v�'r��f��2�&q���T�'͕X����9|�Jc(���"���.f��.�4��S|���C�C6�m?���>k�T=~;��Xx#`r�u���B��G�UV��0}:&K8?��N�q�$>h��ͨt�nW@�����i"�i�A�w�7�"���ȰJY�+�qͨϡ����������/�&�5-�k�k#�R�)J��3j�*�����M<��鈱Β72FC!O�I�bwJ`8�_���+�9����R��k�I+�=-9X�:��L���������震��;V��J����f��gKX��&}��k��_� :}�s�'L��p"2f�?ä���2J`��,�a���}��MɰR3ߨ'CJ������|d��E4�A�ErlJn�ï���0b<�T�R��\�yKa ��U����0�P	!�yP[Y�� 뱨+y����oT����$q`*�f=�M�r�����l�%Ёs)���ޛ�=�LZl�8h2ڕ����	>����y~�	U6���
��^/�xAk�� HVi��k�(�]R9(Q̃d�YnĞ�ш�~�8�&XuL�v��!�H��W�u��A��:ST2���-�>�s���{}[�}��-Bpt�XT�%��?-=*��;'Է��C�*�@f�R������\�ۨԻ�緲�ʑ�D�+J�^VL~�c0>��bSc��&��?N��p$mU�M�a�.Ww���Z~]�r�|F�{���?Q:d�ݮ�]��4/k��g8����ɕ$F�
PQeub6��>�3b��m'� ���yҰ[���H����ף|~�+2��ߟ���j0�,��OV�쪧Ȇ	����R�ƷB K��c���c�B�#'�7�ۿ�����:^�f&�z~�gxZ��9[��\"�$�s�&]'���%m{���]%�c��ܚ#\j,x�1=�O4ۆm��~��J���<����۹Z��B܇����Ý<g�����m�n�W@c�M�Ji��$�ڕ4ĳ�Lp�c��G��pt-�*��\�ց)h4�Б!W;E�^s�.m�񌛿���-�|w���8��j�J���V��6\3�(e�-b�
f,�ebAY�sp�Q/�h��AO��b���8�
�D���ح���'��V��S���g�x ���	#e9&YkP���S/�p���y��?���Ө>���o�]�] *<�|�0�8�nAK4b�6����S��  3���+ �)	7�v�P�E���п�K������{NJ%:��ˣk?^Ԟ<�b����S5c@�K�Ϙ1�^�-ރ�u��$�1?����ඦEߦ���8"�����IW��t�y�eɷ����U^]�G9hqrG�Q��CӦ�o�ȴ���P��d�I^ь-J�Z�+\tA��'�������&��@��
���D ��j5��tp�dmf�i�b��e�����X���lj�CW�֨��l o�2E�B��S5$uQa���XL�Ws�{��E��e��i��?��ܳ��4Z:c�M�k�-z�T�F�q���&��ݥڗ�+�ѿ�FHڣ]���\�L�4���nз���[H��(��0�bB樠ča9Y<.�ty��܏[�������I@����Eq~�1.0W%UI�����X>����#
<X^�4�q>�KH�ۈ,u|�	DnA�]L� ~_����P��%��*�@���[iwb�H�3MmwZ�Ӽ���B�׃<�6��d��xW���������g��}H<9x[�F9����ڕ�{�UHG.��H��/��gaH�R�ݑ�����~6Hp
;�N�V����-�ֳ�E�+�����,��/x�6GZ;�ә����le��z�P���
�5ЭC���
��%[����Lz��(\�o!2(<��4d� oX����V��ө듓��`�އ{�e�n�����@|}l<N~���z���.��S߱T!�
G恖Ijc%��#�? ���)q��	�&zܦݎCDO�UaK�}+@���f�a �91���j�������P�[�����_g�Y<�-$�j���LO��.���Fy
3�t���}�D�5�L0��̺H��:�8�x7F�V�w���~�s��=�8C�u��0V9��eſ�{7r������ە Z��3ٔH�F��cߍ�y3D"�p���wP=����P�Y���h�~ō覲��Qy�))l 'Ä�S���̓��0�ܷ��wo��J��R�`�����b����"|��5�@������أr�'�#k���WC�ǲ��sV�P�s@m��Yf�<�_�M���m"q����-�D�r��ivh�;<�v�y��0Q<�����F%�����E��߲g��x�َb[LW���f�p����*^3����g�%�wd��8���K�r��F�{x��~c~~?��%�|ZT�0v�[�})�'�EՌ�[�7��B<*b5ʐS��,���y��!���L/˰��������$bST`��S�gA�Ĵ���mQ�		 ��+�|V�.���
촋�e��os,�/�	�X(�@��P�ɦĞ
��H��c��3�����l"�g'`�>´��kU���5������_n*{�Eѐl֭��$W׺��[=����H ����Є`p<�ɞWg���
�.���e���B�>A�9�<m�)EŨaS�V N9oq�x2$���[��I3*I�{5�evM;������K`�RB΁~� 7�µB��f��D�������'sɺ�V��mA�$��D�,���ӫkt�<�mp^��iU�p�ŵK��#z��\�ݮ[KS�/r���L�5M��;�om����՚�a}���w�p�h'I#4?^�с=�c����}-J��Z�|�oj�@����\&�V5���:���2�>S��ꞋQ�厭zm��D	���`��s��{!�DDr�-?�{�u��P�V ��L��jD\T_J�{8�U�FDZO�"lj�|�20ѳO+3w�5��OƌܤY�8� ����B�r��o���H"â�iYy�>Y�XLi���_(���ƪ�0��yV�s-�8@M���0�c��pl�eN��%߸��Y~�3��K>��G��z/�%�0�����#�f2�7�2''����=(�:���_�j���42,Ҥ�+��3���k�$ؘq[�Ү�H���L�G��]s=�|�"���֩����iɽF�3Cb�)aF׸�i:�/��=Y��'�B�K7��u�����'_roP�r$5�Hs�v�f]������D�UB�>���0�h2���*�	,ކ��r.��u��î�瓸�B�]�w	`�>K��i�ZL�ْd2��;�s&�}}>_ny��RJ�j�~�7.�S9��´(e�}|UH�	@��WZG<mL|�Qj�Z�zvt��H�E�*(��bW�Ř�e�+�D�0���XՇ`�Y�[���b7͇���ja̹��s��C�0=��m�����Hb�W1�|�yC	��P�L�h����i&[�dV�MF�-r'�0ڴ���d�"y7��9�	��t���^ �UR7�3e�w/�\���+��a��^�)�|y�̵��94�4y.��Q��!o߉�������ս��A$%�Ә����G�G)�j�A�3�Yuu�x�dU!/%���.��GjK+����:�N��R ����