XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ā�u�`��Q���\��R��*缠>��y�rN&
�VO�o	�r��G@��I�I����uES�̕y��q��6��$���
����
�}�X^p���h��d�	ޞ(?]��ˮA�Ҙ�g�c$9�W�fw�ػ��"�I�M�X0	��Q�0��!j�o�Ɣ�>�L��yc��qTƯ1ċ/Wb~l@@�E�����8�V_FIe��Ƴ���������8^8���� �tv�H�vO�����z��o*�+fgyև��Ӥe9b={2�u�9�E�qo��{��h�CU8�� 	p�!����\���~q n��Υ�D���ƺ���%�>���[�?7q���O8vO��>c��ݩ�n�en,�=�n�Pͣ���+ǀW��u\R����~q�"��p7t��#}#��`�*��*;�UB���[�dHi#����	&d"';���~8�X�S0��Jcqz:�CG2VzQn�2l{>�c�0g��o�R&X�aC۪˙�j�.�؃Jr�w��4�Rכ�MҤ$�H�ت�L��"����4�J�[�>M�kb��g�6 1��j�5���R��r��M�<L�'=�Ŝ4�?!`��zÆ���г��?�v97���	��f��{�3�_�������0���g� +0bR��y~�NT�7	d�"s�	��7W�$�Η|�e��J�����G �<�)���"�X���E������o`r?m0����U
��O����__�v1Oy�F$-�)&}XlxVHYEB    10e2     780��;kz�cOB��.�~YM��JNP�ڔISg�A�E��Ǌ��W�\�oJ�abV��2�.̪��Q���\Ҡ��i?n����
4y������}]U�vޥ�v��@���5�j����/pl�	k2�0n󶛔	T�o�@�l���(:�����P�H{��:G�)�q�Ɍ�"�~����=�O��}��b�{k�<���j���U'=8��k�:�8����|����c<G
���I|��7�ةc�/.�t�,���솊KV��Rg�U�p��������\܂�	�R_���1�
�L��#�&wB�`{�$��鞮Dɪ��N�@1�r�?*����]`�n����+���'�`�F��ԯ�Qc�����y��6=�?��r�k�(���~<n~̋u���!���zV�%Y_�4ފ2����1��r�Z�rٮ��J˜/?|+��2r|j.=,w��ϵt�M�PR���O�GY���!%/�D`�����l_��	�!�v�M� f����vT�vW���O�ͫq��7�Z�p*���o�ن���`���,FC�zu�z�
��y�i�4�J�Ie9�S�J�4��tT���z�Ώ0�L��>�A�y�R�q��D�p����\
������n�}ke:�& ���8}>ޥ��d�1� zЩ�2�O���<�o�90�
([����u�h'�$]Q+���Qmw\WS�	�n�r������ҧ%�-�E'{��*�Cس�$ACU���X�$x�J�b���\�͋D��4��Q�X,�Ε����dr�A�7�(��#d��U��qcܑ7&���h"$KCҗx_��]��a�ί^�U8��&:��oǵ�i��fJ���V��(���r'�q�P0W߬�=��{�Tud- ��_IP��aaa����,���1܅Π��A�����צ���H�n��
 ��3?�h:�ͷ�?[���}��ڨ�j\��'��c�A*�����f	�x;�~ �����ɹ�p��&:�b�ц��[��D�R\����Ԭn!Vn���v���j��ъ{� ��� ��̆!�W�d0���'S
�q����==bF�׎���o]��S��P&S�5�q�YHy[��s�6����o��)��y�+ݯӅkY�ǐB����Ȯ�3��1��,3>&;�����y�a�#�����QM�C��13:o�/���C�O�����o͢��>�ʤC2���ee��B���ݗ�8�g�lls����&��Q]LK'�Wl:Wu���1�#6b�p[��hyō�52��BҢB;v���G��s���p�o���}�!~��I�ohҺ&Wm+i�Y5�ˉ�k�����ܣP'J�#ބ߉�5BQ˙�kߢ-��[zV��M707�Pؿ��A���֫n0uo$:�<�
܁r�����w�n嬱�'�_����3�Z�����zf�tؾ(�Q���#�q�2��Z����Щ�3������71wyR�J�4��R��a.�� �:�c?��'(Hk�+e/C4ܯ��{�e'������ʪ���\������h%	ߊa� �^ԕ!4d2�����|
շ���C���Xy�����rH���?V�kΆ0����u��_�=��a�L�e7i��	�jL6�0�o �训g!*xP��/%�ph��Q9;s����$��� �3�&�I��1E��3H��F4���֑v���6�f�2�"��?'x�29�0�>H±_�����6M�Ԏ#��T�T�w}�_)@.�eK9���E6Z+^h~���`өlVȦ�B��j������n�Lj����w�ǧ�PN�	���%л����M�� \3�NL0��=6����Lպ��V=m�"�m����