XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S;Y�D`}�vB����� ��"*K���y�e�	5��5�D@�����������	2�u/�H��#����(��̲�k�����Q�p����4\�"^�P�Ag+	��=���:�q��m�g�>��U�%h�g)~�[����A�F����ش�x��fC���C�n�&|��x
v0z�?^>W���2���5�<���HiW�>��H�t�Ka� �(�
ѫ��Gs�yu��M�N����R���Br��a�ŖV`�z�1В��Tzp��|9�]��1�A��g@��DP����ʟk�g�N�}9	|��׈�Ѣ�ㆫ/CFiGNM��e�4Uc�֤�O�ì�ِȢ���t"�G����e�ݏɒ�鮤2��{B̎�D{j|	���a�i������<����5	��҄{fϒ���]�1��VǾ�[[n
�F��/��Jɫ/Ѻ<� F��;Ш�_�-뉮��a�����F�$��1*�h��F�����`��L����L�GL餔��+X���(y?�)�ߒ�	�{��&8�{ްڤq�y�����J�Xr��-�1����i��#�il����Tl�&�~����ȋ ��m%r�T݉�����9���8g��7�n�ܢ/{*���)�Y�*$Q�e>n:�W�B�b���v��œ�9�a�ia<zK#�UTt(�&N�
��ؔ�Au`JHGiɽ�x�ʸ����{�S|+/er����ѱm7��c��?r"�a�GXlxVHYEB    38c2     fa0Iisp�M�p�A"�_�Iʻ�Y�=>kDHp~	-
�ih��K�E�ׂU�F�7ΜL5F7�r[�g%����^�ޥr��oA~����|�=�,I��L�kE�&��e]��Y��ZMZf�V��fG�$�
����#����{y��4S)123� W+��te(`���@�?�2�#B�_��>�=�ll�P�j��b�
�	�!�'"�O����d���[B� r�{��ه�/.�Ӿ�V5%ŋVQ`�O�0P���<��뀗��w��\����pP;���6�3*��A�\vɫ��{s�ƅ�9�5ڧh����=��m@.?��wLG2qͶ.d�����U�����y ������&#X��c��B����~@��
���"��h���?�NV��59�=��Y%�bY��$�L�Gd1�G�I붏�[�p*r���9�u**;"�H"UU�3$�Ls�@��s6صy�=N��I��]ު�?��j��H������_�������j�6���#AU�F�o�����\�M�:~S����D9�k٪| ��fz�̕�C���s_J��Fe~ r�x���}���b�=��𨭸�eX����"9�~�L^Q;����'���q�D���B�J��6,S���zp��|�F�ga�/'���)��^ou����sV���h����ϛ��^�k��������H4�3zi��2��`�WVk|�&wS>8�h��+-M�� ����
U�*�Q3��r����F��˭mml��e�)���=���(E�7u(��߸0U���C��k�I�œ��;u��m#�:d  4j%��4u�<���SN5�%W��Z�VZ����0x�a��0m�����{��ı��t���C�"vTN�E�Q�`��ْ�cKkô�ܕ0/���©H�rƬ�:��h9�8��[���}#W? tJRC�%T���<Ϗ�%R�S��mΊ����8�Vi+�iscYQ�
���x)��'���N�������S�VS?��g���8��}�.2Z]�lV��;fK�zS@� 
9j�����iv�?E�$���%�0�}�q��.C�=牤e[uA�xp`q6UN�G�ms�>�_���z�����Qz%�GY:`I�6aXS3�<쬀`��<�Q�7%����s$��*GW�`|�(�n���n��V�W�8h+r�z�p�M`� �[Z	�Q�\i��)Bq�J���c]#�eK��/K��I�4���¾}�s��t˱.��Ù��m(�)�˓i芑���
g�̜Bw�M������?=�B�f�v�״��10Y��W%�P���M���E]ֻӫ�w�}����|�,���a4���'��0�/d��#�#ы��#}�bt�}�aC��H�U��˭�I��I��zYdq�/�?�K�+a~���c��2��G$�$]�͌�W	I�ʴn9ϊ[vR9����I[w��Y7,�y����C�V���ӝZ�Tc��ԥY��fe��j��j��J'����V�L�b(mb6Fˆ��>p#XEp�ۇ=l{G��,����C�i��y�d�C6X\,u(�L�V����a=!YO@�M@��\�>������z|������w��5�"�{��1���~�.3�z0�>h/����|�A�b���ם�cq2n�Z�,�������5
*�
�3�H%�M���5b��� F�ف r���^A(I�&��e�����$�wD��,/&j��%_F%a�=�g�����?��:���u<Li2��8n�W�r�n�F��G�}#��Eu\eY���rkU���1s��U�Ϯc�X�ʣv�(}�}q�9v{K�����!g��1V��m��\���:�t�:ts$B�hu=L}����f�G|��� ���f.l�3[z�.�c�5Ȟ
'���,�+�:}��U���� ����W�j+�S��K��������wH�Գ�o��H����Ki�/���>�Ζ(/�	��C�G�bCSo�f�^by�X���}?�?���UM�?�E{�!� �$��������8���	��˛];�A��N��-�e���b�E���������~;�HH���ٛ�,��n�w������:j�I�L�:F�,��`0.��Xa�]��/�.��>9#m�~�t�ԫ��K�B����7���RX5��4�;P:���)���70����U�Ve}8�J���-�@ժ����$)q�?�D�x{��ýIa�̇���f,�aٛ0?��di,��Ԋ�9�v��|=�_5N���Fc���>�<��o8k,֞6zyF�V�l�C|a��׊,���W��}"k��[�2)�y��r�ϖ��0F����8 n�ѳ��\D�jJ�������!gbhJ���֓��Qc/�	���1�Z�	�E�daK�8?@7}]��)6O�I�hv���	,ɥ5��wi�)+�6���<)�t����M���m*�Ges"E��}
U�)R�&j�bC
�%��M�\}��:.��lYf�g�?G�/
��x�D�Ǝ��l�!w��7���K�M6l�ڕ�^��?�Ƙ����V�W8{,ў��d�r�Z"�%I�2�����ޔ���2����4=�-��B��,_^Ͱ�ژ|L~\]�?8��>�.�]�<�D�d�6_3��1n;YOդ1���K�#���P&���:|�n �}RQ}���LP�!/k���(��p�^1�3)A�V��RǎyD�Fm�fF"�Y*0�>�ߺ|�ѓ��Z��q��Ѵ� ���������4�U�������gO��ʶn���/�3�����1�z�Ֆ�w=j'��n"�$�y��3P(})�p�x�_r0tw}Ŗ80��k5��9Z)o��ұ�<K���봏�WQ⩖ޗ���&6=_�҆�o�. ��h���b�Xu��@ﱯ�Ҋ�Q�~�%g�4� ���ُ�{j�Ga�txK�1��a�<�鍈������so��-nu��i��*��Q�k���J����,����h+G�h���y�����
6�D(x@0�z����^M�q��V�#�׋�o�h�Ө�����}�j�<"�g�t�D����_�������K�#W�6�T�J�/���8м8�����U��¶,��N$O�):���ҷ�L���7k����#齇]%��˷M�_���U8���j�<v(Z薾���V��G�"�����.覰*%�>u��e$b�_��Ϲk!o�� �&���^�L��L�-XpK{(�M�`ү�~�7�2X�,�[3�=S�"{�
7�\=v��G"�w�jc�)=�à��[�@�� �J/��O��$����=g��qH����q��eB��v,�
ܴƱ�q��㸳%����+�R�f�K0c�6��w%���U9w�F8@�,��7�@����t����'R�^����?O��� ������(`�X��������<�Kx�z���)?2q�}`V�,5����&�YI s6Q=ŵiq�>�U���oW�P�ߚ@;�b½V�����@[$�ڂԨS7u.�A0|�<�)?����̰�6V�z��49\0h�d��jS�{�lG	�y�z���oS'R��\Z<S@�d�+cƖ��%�ߍ�r�2%�#P~�F���QP�A�[Čq/}б�uS*<�ӽ2�}D7/�^�j�4���,�WQ[q7}s�HD��$�~��� V2�8�ڮll;w���Z�W��lf骕�y�p������~0��/r�g����rY�2�;>�J ���غ����gE^eZ9��*[)__��9�L�-*�o]�m�ܳ���F'l���ڷ6��CV^(qg7=,����o�-�`��Ksq;â�N�"�>�p%�q���F�u��w%R�-��d�.78