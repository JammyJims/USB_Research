XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D��A��ےT+�ȷ�+u$�[z�.hB f`�GO�]>Q>ɸ䋿qq��F~�$"E)�si�y�Ry9	e[WG��

��2L���F��R*ه\{D��  ���}|���@L��1��@�mSV�`?Gq Q.�ϕ�����ˇ��H5����2=e�⫩fce&E�Tn����q�=�ʶ	\�l���r�j�_�d�i�Q���P8��3�0'@�#���J��b�|mz�9�4۵��]��ÔϤC1/|��O���)}��-���b=�5��Fs�ZY?��B�7�\!��"��l��'�`g����Q�
����D~<xg\
ljr���ֻaI�6�*�������0��Z L�^�nb0���,��G�.^���_q��( �nt`?[������ң�G�Z;4���zHD�v���T��F�ro��v���0t:�&w��4ܣr1۫�ǉ����#��Yr�e���N�Rq��?����	Q���_��y����|M��2��_�T��q4���bd��S?_[y'FuY�_z����_~F�b���֘QyxW[_��Ɉ=_&!�L�S�n�`�8�X|�4��x:�I���7ՒP����:�����B��N�.��P����M��3Eq�`!&E�n7��5����,�v	���`G�1b�����Ė����w�g����k��nm����rڷ�u�#i�ȧ,J���Qc��{����M>�M?kGٚ����z�X3$��lأ����.��*eἀ��moʹoXlxVHYEB    124a     780i��ɏ6>u2��>�0���GZ�J�V�g���)�xs�0��b{�"9�Q[��ʁ��ޛ��]/�Y��;����bF��!Y�b{K��I��pE��#u�����A�����O��7*�a�|�WؘC���D3w��٭�kiB�w���wb�Hm��I��n~@.g��`����M���:h����'a�b�L��n2�;+�S"�O��V��]���O�L�,uu����i>1K��pj,P��>zEoC�d����������Bn��fͪ�Np�!$�m�\��Ą�R#�=��)���oYl�;v=x���/�<�C081�B�9��za?���R
�{���Y6��Hmғ�j�\��,��ʯ��X4_w\�hպ�)5�݉e���b�)�m)9o�M���i'�{�5-��7AJ� �T^�H�J�H�w�!���2�wG����8L'8�r��@S�c��k5�S�;G��+� F�.���{{����8O'VǨ�d�ꦨ���Q�<�U�sM�u��T���{-�FX�/ǗYQ���5%�&���X(Du�Q�7��%�[Q"�[�'ݱ��6�����3����w�z;w�H�F=ib�L z$�;�7��s�i@��m}����z�~��ҩ��s��}7\�$"��D��q�8(�Ӗ�d��#^z��2oq�A���㹘'g� k�XU@���}��%�=$��E̝�H՝oG$غ?�L&A�#�=�S��0wc��n�ΝcQGLi@O�O<]���h�ptί�dj��M2S�z/����8/ ��z�>���\0�0Ƴn!������1�wЕ�ߡ���Ȫ&��	�q(kUE�����>�L���o/����ޱ3�!~߆���u�p�8�6?�5�ro;j	�󲁎�s��)�_�\�U�N���m�Ry�������x�^�R�+g�Ǫ��#��j͑�m¤�L��w���97��Z>""@)9)	��r�2w�V'��A8�0��ߙ����w�<�>}���ر�����p�c�#��*'2 ���Ty�p�92�w�*���Z�{��A*H'�G��K0Y�A�9���pt+���6A 80�B��WC!�1,zv��-2h�癸-�Cע����<3�J���ĳr�ڨl#�4�oZ)�%H�)}�����g�[`�0n��̕>�w��i��A�?q*y��{C�OĞ��p�O�+�/���i;8x��>a{L{����b�mޑ$o@=U��{�x=���8�Aw���E&�����QC-�V�������x����Zx�أ��
l�������[������4���{��?ޑ<��G��6�q&��>�����p��+zv�����@�l��!�Ȩ��W\n����ÚY@H�!=��\����0҄m3��;X���S����lm5���>��,��A��Hmx� ��%GQ�#�S�A/H(��88kW�|rv�nh�Z�7p�/�|l�_��GY�'���/Gxc<b#�%"�;[	(�?(��Ѹ�/b�;q�B�I��k*��=`vy��ڈJ���a<�.8�F���@x�P�f��k�$��-��5!U�����[�Q��� j���Αd�<]���2��8�O'^�C�i^�Kw�@ғ@�~1(.R�*|�Z4�	�@cA�V'������~x�\x!ꎦϔ1��\�����.���}��'��+�d���i��aL'�P��!��t��lx�(�����������������w����'�P͘Y����TjT*2\���?n�֓����Q���O���Ǒ �8�f�C�?Ş<�sw-��E���%m�Z����1�/ȇPB�(���gU`,���	���y��/��B2�3�ŋ[�֡��%�