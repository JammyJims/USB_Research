XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����w��S1M
�H��+�]�*���7�d��3��X0<�S�Є��V�ٕ%:W�@��B�2��������ۢH;�e�Ҙ8^�K�N�k��B���آ_��Ҥ��L-�0�"�HBv��yy)j��.��o�@k��6�P"6\&2@�s�8v.��|����lG�κj��M�u
����2u�`�?|�VH���P��O�K�֠cz}�p;�H���E�ʯϒg��ҵ�R$C��S�����c1`(߆�t�0-�I���"��DL]İ��NOn||��F�
��������IX��`��1����~��m)�li�$1Z�9�E�ZϮ�1�.!Hf_�>���ťzY�d=T�J-��{� ���3�	����s��\�<�&���W��' ��ͽ�4�ا;��r_'�tņ[�Q�T<v���\�ƾE8�!n������8&;x���O�RaB«�0�W�)M�)(�ăX6h���1���IO��z
Ƴ[)�Y�8�[N�����������c��?�޴���ԟL�/���yR�RY�)��*��q�'���gl�;����ZY�h��N��j\~KXМ�:��A�̏��%*�Y�^i�����a-�lߵ��F�w8ɒ����ߤ�P���X,9���7��>k)�A�"#������'z^Pyр8b,��Q�X$m%��U��$Zr\3���� $��]�� �Nw"�d�n�����tꡉ�9)��s��V����u)˨c�/�<]%&�m���T���K�X�NXlxVHYEB    d410    23d0��X#��5��Ծ	F(>ܖ'`Ä%�sx����w���АSwa�3A���A&cj/Xf�6V�0��e�Er:�ȋ/
�� ���U��ᑫ4,A����o���l>��ґ��W�PM�	����f��_�{�>��p3�IE�fI��$q&�H�/7'�Ut�H�"���T[5�~���ޠJ�hF����@�!���ZR&-~k��,f�h��a�U��5��e��gJ�_>T�^/���n�ꐱg�W��|�OL%������4�dx�z������o1�٩5��:�x(�ҁr��+�*!77��E���Ql&�2_�Tsh���-�v<P3��м��;g��VX.��y�/��;8�����r�S��rRV{�\�EƋW���O��^ee'6~k-���sYW��b�w-�(��b��#�g����D��tފU�T�oh����P�`'����|e�E�y[geB�G��{�1���s�!�����6���XĚ�^�\�q�^�e�PĄK�/���/�z��»����<�UE�9�`��?�a�z�T:�	������!�K�)��/�F�ˁ�����lu~�k�{A�����)+F�D�_=6����/��k��S%�7c���mL� 4�t�o.���v6��:����}��Y_`�!��Hk�5B6�j�`-�!y�d�&xB]-��z�������(���FN5�fHEԏkFI�WFn�!��<�M�P�m�Y�u�zN�W�6r/;��Zu,!�~{�`�ڔ��m�l}r�wQ��P"<Wϓ�Z����P0���g]���0���̸��o�{J<ؤ��N��tE�!À�^�VYD����S!���:b�q{R���^����R�ᗙ�'�m�w�+cMfh��;���s��[�ą��}ү$O�'�3�́�r$)��e�����~l�ħU������疼>ϐzwO��S9��ш.HS|YM��+��Z�؛��%?OQ��`��|D���'|z��L�^�7���� ��c*��q���բ/ۈ�H61�����I�~P��>�B�2Maѽv�'�ߙKХ��Y<��qa|�z��\�� ܸ_xUH=] �j�����Y���XkU��.=!��$v��5�(��6Kj�.B�yĤ6��I��E𗨬�e2�iS�F#`��R�(ē��?�_�"�s��h)�c����WC�+�d���EU6��^�&Tz��~��m��J�/ĝ(�!r!'�]}zms�m/��	�4�/0����- 9e,	=G�	��*�:C��t��QdfU��R���g��h7�e�j]�FݜqD��c~��rf;9���`AU�X��R�J��d��y���8pySN�I��H�/&�R�#c�����:0��?c�]ΐ�T/� /ی0{3���� �Ƚe��cɻ�=j1b��]���(D�Ԓ�VlS���7%�!��X؈+k����vCt�!��i�2�j��"v��hq�I��⌔�d�+]�N�E}�h	!ʆr� �2tJ@HI���$��x1iDFaV(&��J��ڞ%�k�#���&K�.&�{��M�F�zs�(_�o�)@p�Zn�
6�er�V�	��nxvD����c�@�#�!�n��]��B�B1�}�� ��ge���PV�'*�Z���W�"=�O�Clȅ�#4��5�l�1���eoZ�����=�7-�R�9��'�c��%3��5��Y���x�2z������{���;����izf��B��ʶ��5��rE_��Qoh�/�^�,���k@�N��E�P%w|��u��Ş��Ր�{-�6�N�����)���F�������}>OX�c�%~�
^�5�CD��<�3�8�Q�7�p
h���įZ��Ɯ�:�+�(D��)]���%/{��ݖH�]5�d&��Kj�QY!�`�3Q!`Ĳ�k'T�<�+ooW��đ�v_�� ��J��h:�Fjǿ�
cgk�A'E�#�MP�iud���H8�7�U:�D;#ˬ2�6I�֔@�K��G�o���"�h�rf��H�^�����(�r�\u�����B��Uje`cmSp]�e(A���!pa�Dƾ��XC�Tc��E��E�O�F�f�ڴ�)c����&#��<[Ίa��A��h�0I!8$���"�zK��}�_�l͈���)�T�9)/,�&#���OF�~R[�[�w�>m����}��@bh�q�:f���������2�=�,(ţ=��ɘ�j+x9='�dHk�F�mʧ���;��l�sc=��h�_��e�c�NfK5��|�%��\��i@1*/?�P:�6�I����cd���m�$�eO�Ë�3����u$�����vߑ]��k��ܴ�A�
�Q�EN��%2~�@�n����1"�O}�ᛲ�~ �̶Z>�s����K��6�<�l�qj�8���^Yk�)F7:޿h�i�x(�3�,l�B��5��5/��[-�ox�e��	iQ��P|��L�/����f:>�}+��S�Ї�w�B������T��l�h�Vo��_�a�q_��FÆA�T�~�9��)�]����1H�Jvm
үo6��#T�m(��Qq�i���f$�j,f ����8��d�sx�e[���i�I�NS��/��һ5w��8���a���^�~;�J���W��p����\��64�.�/ى�2���+ؗ��xN�;w��n���f��#!p�x�y��W������q�._�c�����ehD�����[?���G����s%	酢�4K9`�%�N�G_w�H8ٷ���㗒Z=����cl�<Ay��e��~%�!_��Nyb�?�$l��Bl���wa��-���0�F<H�Mk����P���R"ҭ $#!
bɎ�j���֝pƘF��?��!�����]���v�����So�͇�b�$ּ@�0T����]1��*�*m�U������$��������f.������_��nzK	���w�?��(���ʒoC3�mu|�� ���h^/�aȞ)4��E3[��D�5g�'D���%Js/�oP�\���-I��Q���w3Y�W��q��uCp����8�C��X�����fI�c���	0��*�F�6z��3wg��OY$��7�O��\�]?��n�hb�y���U Oݿ#|�W�<�O\��H/����)#�&��9�۳�y���(t�!L��8����ڂ�U�)�xhz<�g��(�;*!	�n��/Օ�5l�F�i��?�$}��$mO��"Y�}m�va!Y8;0��r˴;���e��4DAH��f���^<5�;GU��x��
�3��0
��?�����#V��6�3���h�#˦i�Z����%�?nHH������o�luC������NL�:�YSLtHw�F)��B��D/�?�e��_Z*xt����Rw��pa��pB5ߙ���D�a{�-���5;��$�(-�ǁ�+��^�\yZi�Č���`@ee�P*��� ����iSWX�@D&�)3�L�k�{���%y� 2%����;B(�H��s>�ԙ3XI��f�V���FҐX�JBNB�(����3êlB�4$��N�+����uY��$b���N���/�p����Ԭ�;�yt�YnH.�3��ҭ�&�Ŷ�Aa�筅�[�B���Ǧ����L@���8�H��tk|���&(j�n⫨eӫ��=�G߳���Gy����(��'�<A�S�cU�z4�"���aq@a�&��c~v�B%����)󼦚���,O�[�\�pf�o�!7]�Q��>���/�̺+^�R�R��h�z,�P��l#,�D�ď���:�S߬J�i�wQ�^+���~��wc��1^�+�SZ6������~�����q�ݐ����耺�2�o��k�L���t��!��Tq��
CBj�I}ژ�̱��E2��b���y��޼?Fv����X��{U����!�.S�L
�)�s���sPB �㫈s �����6�n�A��G���d�P:�"������#o+R��� ��,*����?$�Qo�@�Zts���O� �tl������a � 6�d�ߔ���{=<��9K��,����V�E��3c�ܐ�ڔ ��S��jCE!F�x��J)E"��T%oC��fR@Lh}{f��
����Kv���?B{��b� ��ޟ0�]�И�x ��N�k�Y��?
�s��J���[�S��}�
���о�U��`5�t��@����*��Kh�?�ٮm�'��3�#K�ۈ�����nİ����
������}�]�㛜��Б1�qV�|	�b.��H��D��i.EϮ�)oR���IIw�Ib�K_��0���iH��!�m%gx~Oޅ���,0�x�x����}Z��,y�bAx�Q��&I�kS���Ñߌr��IC�%Ӭ5]���OBI�;'(zZ�s��g�ڏ��o�_Mx��JBL���ۼ���f�^�Jt�U	�SϿ8?�<1�1{��2�s�%�,����3b�L�C�H���W�L�y�,_ѨQCh%����(�"���G��s �쌌<O��9�F܃� ���H��}[)&�|	Ͼ�x��|v�P�Di�U=}wB�!ᱢ�h�i#����G��)��z��K�g �.�r���L;`�3�r���I���*��(��!b*��� *�~�����e��g��]��� �q���k��i��rA��N/�h2��|:yJ!�HY�ą���cxїn�[�<���YL"_�ѣ�sP�A[LGg�xń�.4���T��Wx��f,A�ǍL �����M�1�����$�����-U�YA *�b��l/�tb��������EĜ"����1�{dQ�@��c1�<9Q�E��'Z�tS��w��#9E��he� jw�y�jRL}^���nN�͂�� O%x�Tyu7��v�Ѧ��Qb:������5���D�5G���Å�2(�T����&�z��,a��`mkKX��L�%���Pwj	uN� H'����4|Jhr�V#�`����,jrV��QB� .��j�ԛ�Kzp�Ć�������͢ �~9�"V��
�r�~_W���#`԰��>�/[�sJ�� nSn6�Pu���V�WC���ͽ���>��;^G L5�� ��3@��N6o�G,�����K�����!�v�:�mDxr�a��o��zK�t�ʗ�V�]��W���p��h<V���'ς���@��kMoQ�iH6����(�h�j�<Y�|j�_��2�y@�N�e.(�2�񑑏.��/�H�.�l��=�&��<�V��`U��S{#�L$ɋ���x��QI�W�k�& �RǏvRi���N�f�x��B������lŌ�N��W�b4�����T�I���QE�� �J$��j�{�g�y�0,��\N�|���1�ͣ��SYX��9R��	h�Z�q�VH�����t�yD�����Ca%��f@K��p������@ĉc��h�V��NFTu��A��LM�d&\�! ���x�ˣ��L���ۯɲ=J�ߨTs��+
= ��.�͌��S2s��/�eAy��Qѳ0�y��s4��F�����gy� ��f4�����A�}�3�c����*��wr�V�_>��MnEE�(?D��L��56|��E�hZd�,��npi
��y�O��[OΫ�\i�*���m|�����Ǽ z��8��	ҵؖ���E��#�w� �� 1��2�%��{�Gץ��� �C�������=p`翷��T���:��M̗+	���~�N�R �P��qJ��d��%���XA�n;^����Q�58MrS@GQȧش�B��Q��1S�~Y%C{��[���w�>��C��(�-�s�*�4:����H?/#.�q�uR։2���2�AMV+�.%اl;3����^�=0#��kΐ��r� �9���ܺz�7��Lp�v9�'q���*+&"k+Z�^�q_{���^υ	sࣃT�2o�J��0K�j2��^�#���.��L%�h�^(L�;����%5��}�(�q�
+�R0�,���Oq����\�+}�[�N%�3�v�׼�Z�wX��(�OlLr��F ��Olڹgx�����po�µo�'����Bxvvz��}���ҧ-y����R���V2���K��Aʹo2�4�ծ�k��'��b`̐���E�^j�2��%u�������PQ��2�����p!F�8_���V.!�DuD4�������ǿ03U�Ӫ���ۉب�m��U�Q+,����\�m�nn��	BC|�+��3X��`5=F�g��R\�f�핦���D�5կ���I�1��O� ��N���&���юZH3T��Ԅ{�&ᴒVk0#9���G�~[��Uyr�6�=��S�M�U���ӊ|���ݰc�d�@$�JG�U���� I,��0�����"�"�ԟ,�鶸��^�AQ���c2�"�S^�H��w��
x�,hɟy��U��Q�" ^���7��QO�t�C*�FG�>H=��u��k^'��W� �����B����� <���f�u��E�)ֲ��>�s�Yr'VS�nS0%�����0p(q%݃E`��L��>��<��p�<"�T�p��$�
̀Vz��Yn&���iTܽ$�r��|�)��@�ys=M��c\Rz_e��}m�&.�T���"G��Op�Q�*��g�Hz:���T�s�?TX���;����	�ucQA����H��ǘ{W�i��b���ck�D��j�j�?�`��WD@ԓ�),O\�|��=��[9;�l�tvGL\]�H�^2���ڤ��o�R�e�3A-7G��eܰ<#?z������8�T�P`����@��5����:��Ɗ�Tb8�+s�wtw�WP��o����tه���5\���p�����%������g&[WӮ�.l�(2f�6qF�I�%�Ъ�p�_��5���]0	ү�!Ԫ���7��S1ݷ�졨� ��x��֐�Q�?�����f�;*-<IA��	9@5���.LsGdP�O��z�FqC}�3�Wa��M��4|^+��/x��P�)n�t�uR8�R�=�TfjD�(`�3�n֌�`�N��)���ڜ\ì���pxqj�8h��
-#��;�'4J�h�������!sgCG�.[�D�58:"��k ɶq�= ��!~܌|]�^�������}�6�%W�H����]+3����|9���D��H�l���BNٯO~{E��.����߀uV'<M�h�_�؊_C���9�&�Ϳ�p-۴�r�9vp+��
�ԏ4��:6@�mQ�I[�%�/u}s�X�������,o��"�e��D�Gp<�=���@N���o킂�)�f��YJ�Aԗ���w�K��׊ӏ�:�����G�Ha3�^;Q��������{Uط�r(F�&�`��)��YA����Q��v���r�_�ć�&�9��ס��t>��I�d���Akn�/�E+���v�2�����\K�y�A?YOf�jQ𢡊�^ h�c��;�9��DS��rP$s�@�|�C�EHߑ�}�琞�� �:���D��`���/��Z/��y�e�Kt/_�]�:,N�G/��~��A�d�[R���'f/��ۦ���#XOA �	����ew�A���s�+�_���,d4��y�#\�ť���si�:�*�����"O�@�.b���C�fTC��V��.�^�� 1���MZ
g���
��۽�[�rV�bV��̰j�(G�u���F�o�F�PX[[2H���1I�lE�ʸzθ�U���ȦN�?Q$��k�*�3E�_�kZ�1սVV���@x��6�Q�ui0���3̬�@DݲO<Et+�>��^>G�'�\i�f�щL�AW�¿�[㜀��tu��9��r��51������Gߘ���+�jԳ���>P �/��6s ȡ��&�U�����=��hL
��)����j5\U)i�����s'i>H>�^�d_��QR^�Ό�B0�7E6r�@��תo�6�s�q�o5�;JW,Y�*R�\�u����P[bG�z�I��#�yWX�r�(3�	p�W�%9�|�NC�P���������w�F�y�M	UX�-��=�'ds�>�Tu�T��K��3ј��E*�Y|�ИfZ�'&��"�I�{�{|�a��b�e�.2s�%ew�e�����>�I�q�ݖ޾�ȶv��Y����:��yj�9�3�i�B�<� �촌L1����^��_r�u�[K�Rׇ��껍~6$�QÛ-o����=�nz�WPW4}f�g)MS؅DPZ��E�`�N���*�BL�����KȂ��Mm�NG�]4�v�����)�Nc��h�(��Υ���@�<+���ڈk�qȿM�#�@���+@mm���KS}��{D��[��"�as���M,��ʴ�-����$m���o������2k3���{G'������8ňq]��&:pf
�X�����r���>,������*2F�)|�f�bh6�m�L��,�(�A�6Ɍ��6v^,3���Aw��2�9����ԫ�:�c�N�0��\1�-Pi��A�4}&�+�@T5|O 6�fW�C� �
&�%t��p�,��'�^o�CY�C�tX�*�Jv+�v��b�O׷�y�K���(�^�U����+�ܓ�}�TS���L&����g�R��6�1J(�� 6�vϏ��i�eEyG����,kϫX`¾�{}����>ǰ��66���UC,�.ə��)'�}�SP�8���A��%�ś�ڑ���JK�/�N:S�	���
�n�E�%�bn'���X�˛h�?NQl��o����V@$�H �h�J�.��ڇ�F�����`���A.i������?����2y�;ﶹo�}1GD��y��w��vßB�t��W���aF�����s�&Aa.i�V�[�EWW�a�rF