XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5��9��eF�I��g��������s�#��0�VP�@%u9��t_��I�yW0}o7d�Cre�e��%;2�t:�{}�_DR �O�'I�hf�f���
Hu+Y3Km�>��}G����\͕*���]�CP�����1��T�e�#���(�ЉR��i��%��)��*k� �K���(�����@����R��՘FP�N$�U�����j�@�F���e��!�FE��-�[J���K���B1B�8�=�
1�G���]k��	� n|��.���>A�fCǗ� �K�t�/���庐�¯AH�suF�v��Lѽ��l��i#�ä4$c��
��>齤�x,�5N���"���������`"s����Y��˸�>:�����-Y
:@�A����HFY��&�LU'�o�^�Po�#
h���T�J��.�N�6/�,� 	�%����y�Ƈ������r�i���L3 ���� �p��n=�'uW�f��g�}�j��Az�|~9�	�g����d����R!|e�3Q#@�"�k�����t����~��.���â��2;�,Z�+�4
�l�:�������%��靖�t�p�z�{��h%��K�M
�R�#�˪�ժy�Ph�[f������'��(1�G��m��]�%������O��v�q�EM��1��Z������ $5h2J	�1+����=���f��;n���o#'�z���V�J�7���Y]u�c`�!�,;XlxVHYEB    b17e    2020���7 �,� V�7�j���8-���A�������@����# ���	��ӱ$��_�_'��iQ(���>a��ظ���TѬ�؉E���0x��փ4D%"?Β�ՀQ��������ѽ|��8�8ǭR�T�+2�8�jzmב,#�v��N��!�*"�\ ��NA��T�N���zf�y��-�P<گmn�W�	�[� P�}���3�mI�k���{eTi��w
GD^��9���φ.�*sٚ�_�W�H���y;ﻷV�4�)��7�a���v��bd������w����嬉E���K�xn�G��Yeo�/>�Ӎ��`��o8^�`�R�
sۈ+;��Y刢p�902+��t+����o��y��Y3t��u�/	c���ƨk,P�����9���Zs{wOCc:�~W��U$j������>U/�H��p�k���AЕx��=&~��G�"��p!s|F���g��U� �����^�	&��4a�
0��m�R�>�tOQG�����p���Ƙ�gg�����+�\���A`������_u�t0�^@�Ym,-��AM�ˆ2��]]�9=�ف}l��(~7�+u��6���.b��AcyBe����zF��^r���[c�|fN������3�=�5m���#�Bu ��Սd�ZQ?��<UE�cRx����6��'k*�Y>S�H��Ur� �q�ׯ�T:fCB�HJi94)-%�����u����Zl��r�p$A�����dۗ��0��#!���h�ZOy�녋�a���ՂDi�=7@V٪�Ͻ|�����.M)cj$+��� ����S@��]���lg%�_d����PO��3
��!� �u�����p�j��������숄w�C��o�)K��n�D릚ܠ&v��έa]�'�E�w%��!�3M��_i��E$x�3*ll_5��eR���seX�Qw}j�������@��~z��]1�ꯍ��3�̗�Z��n� *q�B���2W���p�ћJ�o�l�ѽ���{�7S�_i��*}����|��j��LM�����*�����Mb��(�ݑ=�t��3q�1�Z�t8򻼃��~تIK�g�>��u��~�zAdD̥���Z�Ԯ�ލ�ԕh��*Â�]}aK�'B��bo��o�3�5|1�*6��v�
Ok�@�̏z>2���ش��0G�^�~̘���%T��S<�� j.Qݣ��au,n���j�(���U���ޛڋ6��k�d�0,�լ�{����=��@��!Mf?O˂xr�d'�+��A�6���#RU�F�
��u��������x�~O��@lQ��L
3�����.h�˹hj���~W�4���)s�V�!�+�R��p�غ"gH��!�GV�����鲶���%��r�i���`Y ݄FطR��>��Q|Q��[S����Iچǣ;f
4�Eh�,�䳍·��ɋ��"�cyW��jj|p����cD�-}�5�GC�D�{@.X�L��F��g� �\��[Y��Z1Q���h\mDo��B
��n>O7|���ڻ{�K�M��H�B���pgL0�S���\�,s���=�$�[7 [�?��;�d[H(H��`�o�\���i�=@�0?�]B����'�$}FZ�I+��]���OC�������Hr�*i3p�Gf��q�ܽN�����;NM�U=�Q��hӻ`��:�;Fd���-d-}�u��9B�'r|�<d"�z��g�}�?��e0�O�bϐ�S
���!.��͒R@�fbD��ũ΄]���O�gz�ֱ��
�H��.�g�������?��\��)�wUH3�BUeP	2��3[C�����Ƿ宲���m*]�]:J!�zkj�q[�yQN�'�N�% �vWI���t�4D�a�������?�7��!<�.�̻lBa=��	��J��j\��jw���+KQ1�J���ֳ����̀����<��Og�c_�ʈlY��$."rՂ<1��Pe:��i^-�B[��H�g��W=n�Qi1����3�7!9.��ܸ;���O�m|鷛󰸳Ƭ�"Pm�>-����}�������5tҧ�K�M��'�R�i���h'�����ő<U�\Xڈ+F��6�p��Y�XX�[c���.H�w�z�ΔY3h���p-��=&C�o1��r>0��Eq�+`rT��3t�I�.0T���1 ��6�n��X��cfʿ��"�>�x�鉗�E�/:N���wE��k�>�͇��g2S6O��k��^�1&�s�[��ZV$��ֽ�q9����u��6��MxL8�3?�4/�H0���F���NH#B����KS�8�u����@{�MZ���"PGn7:E��ߋ;�Xd��] -G�j��h6Suڭ� �jՌp�w�٧�#�&wd��Fȏ~J�P}�xw�r1��۴���������;�����V(�[$�B�۳��P>���#�0t��9���s�h��π�c�g�Oag�0mWQgL�D&��_Qg�(_5�y�d�ChH��u���}L*�?a_�����y��s�3!Vr��\������a��~��?K%\l4�y����&��)���1�o	0�P���g���Eǻ�&=.���-�������͢$$p���wt%�Z�O����$�:*M�\�������Lkoݒ���ꃒ��|�>��c�*.=ӋG�,��U��RTi���@,1(��G^)
Q*#��t3�5�f���^[]���r�:��cJ&�$��WW��
x�M����M�g9Es;���<�����xx�%�U��W$�G4�����j��X�,g\���o�2n�nG��d����M«S�˩�	��]�0d�̩U?���5|
� �%Ylho�f2J\��h#߱�ދ\���b����)gk��̎�AѾ�Yc�K�M���z���,�r�c D����=�H�v:���=�|�L��?IP������%����{�8@��ˌ#��0P`<, �[�}������Y�V��	�} J�|�$V�CZ&��<������Fݤ����<��w9D
�z�2��O��Ͼ��}�o��W������ճ�o$�ۢ��(w��=d�[Dƌ�
w� 5��4]�j���P����d�$�X���@�8�g��ž�����-�8��]Ho��i"��n�>�O�P6xFV��V�:^p�2�ey��Ox:�t[��n�����Q|.��
���x+��Y�k���*h���b��g�ee>���Bh������.�R��niտh*szj�%V�z��~�����kPU��F�#�cl���*�i������)i��G����<
%�jY5��+�I�hj��*D)����lM������NZ�S�;eL<���5��ݘM�['�7h�P+��D�y�D��Քsi��ƶ*�wMK���ԭ.b�Öц>� �[���|��Y\�H��g-Pz��>���5�Rf��'��H9�W_���4�̰���քN/X5n>�c��<h-�h��<Oi+g~7�9���>�r�o�V���U`P���7S��l�k
~iw�t�����V��y��ýx��l��pQw�9�i\�#.�R�~�2��V�6A��7Ύ=*<�󠈭]wɶ&�=LC�kwċ��#�K:~��aC�=�9�6,zqg��󬥁��a�{}��n��Boo�,�naA�����r�@�
�x��tJ�C�$6���{X��}���:�K`.¶ �`5�O��5M���B�5^|�{x�7�y�W��Y��� (k��S);��Qy:���ϋ��Ԅ�P�7�쌭����"0٦�{�`|��pe�q5A����&T粩�)��1S��*a���r�7�t	&�F�kp]�u��E�����6��Hn��j��}��|+kW+�F����
X`����bZin���)��^�ֽX5�t��*�WTz0w4����(��W}g��Vh�?�$�^5uQDr��H�V�x `z�^X��	_�7�3$�QK�V�4)�d������?�Ҧ�K��k�߶G(O&
^�L"�a4w)����w��D�ë\5�C�h��ʸ-fr@�G�_ز+KY�DD���f$�4̹R�5Ĉ*d|�Kc�!&:&%��g�*n?�����O�Q7n�5��0d�n���1E�Ɂv Uw�+ȱ'Y�/�gL�2�Q3x��<����fYy�t�f[�j!U#��"%��	z�gV���B�)qt��:�I���Z^"����M�ISh82b�d�5y7�^3���&��r�o��Cf�	K.cE��������:�`�2��h�x^�B���B'��a������K�܀���/�ǔ}��
�O��)�{���I��M��q�+����H�L�x7�[b&� �	o&���OiGf�f�s,_��1���>�=^k�G�zD��ny��wv^kD+_��^��z#�#��p >8X�%sM撴�)�{��ȍ�V��1yz5j
JK~���E,�xTf�o�I�ol\P�%I{δ��Y�؂�%|�����Jn���X�C��`�3�m��6�v�W����{hu�(��H%�����OU}��܃Ee�B&�0�?�~w�B���/��W��617�;�I���>����0���,v���3�x��D� ����X�<����<��ȨX�*u~$��b�%�pM}왐���62E�����F��9�-/�nM QW���
A��VMN�@c�S��;�\��α�C�L
}�C�y���y�NSm4$��@0���� ���&:�V�]fc2L��6�ѳgאzy�
����|�����(�������+D�x�}�o��l�"(Oa�v.66A�������<S�g����	�y�lӁ���\��=3v3.����f�^_���lN���(���'~�4}�
�;j����\!$���k�Z�"��3��ŵ�P�S�^Ft�=R^`�O�����쟘�۳-M-M��=������a�Bu�Z=9Ez�oW5���U���,P����L�Ǥg��o���n��YUl���YD�.u�hRȗ��=���I���.&��]JN�7hM�q�K��b�t�}/sK����Y�8�-�l��u��W�@2,�����7����,���C�7)zlu~�΃��_R3)T��tuX�J�����Ο�k��$�
'+���YA��O?�0�)����㱭�cS��x����J�'N�*�t�	�T�����X��#��/�����W��5�8���s6�Q�����hJF{�]��lF�����~3[S�~F�������=B���;=ܲD�pM���$��u5��H�1"�mP�,� 7!�]̋y�� ��,@����XH����o^|�	�9��7�D5�w�lW[(%(A��`�M#�w1��=�Ǭ�1�aj8+�y����`��G{�J��C�V���\��J ����D�!L�|���I��Q�����U����#��e����"̃��d��1y[�R��3�~��:@J��?�|�d�1�J9��~��)3�YXZeb;�lӡ�j V��0��z�7�-!��)V�)]�"Ã0G��7"R���ͶY��hv���ҰH�:b���%��ί󒉺EÈ��uо� �]e�U��v��gQ��]����7�.l�=˸y[�K�]��l�%�:��z(���
�p<�%�z�	YXY��A��Yx�
ʋ�"Ԏ'�j�p_4�
-M9���ڕJy��Eb��h��:H��F���fAr�7[~6�˃:����5��{����j��5S����3�cνTy.\=/d�f7�vc���o��DExt��N��m�a7�f��N�j�d!^d��_�-���U,QA@D��f��R�6��}��u�d��jC�i_��x7����5~�]Z��bx�:�4]76�
�0w׉tm�/<oZ���	]��b�t���Z�`��;s=� ������
9�fO?���4ǖ�1�7ߪ���sԀ�M����ٮK�nE�#(3G09B�W<��x�m�~�6�k;�2!v���sci���ϔ��>_�M��Yg���y���	y�����9鞔�b���8Bt
>��7���ǭ@�{<��jQ׋/r�m����t�^+p���g]Z��N��4l[_Yn��/^&��l����}NIV`9�^�,�K��(��k�V)�c���ԫ<b��z�Z4�>�y���P6v՘��9�B�9���9�]) k-�)�5� ��{43���ϋ^���E0{#��j�Nc�k��es�|f�AN�^�gt����hK5-��B�v"���+~�i�#��#C�zU��faTo#�5�_�%E3W	�v!��������%f� ��l�C
�(w��_9OxNb�)r�0���[�V��߻4ം�!�17�?�.K���CA����o�w��������	�z�����{����8;�e9�n`]�X��3pk���N��v�?��k� 1�-G�F�"���Tπ$�e��07Y4}�{7GFT������[:��1]r�Xr�|��K�F���%':(T'ן�ϘŰP�+��'�ߗ}Պ�L'|������{���r���Q�j�T\�u�h[c	��.�����6���a���yY�b�\i�����*���qů�����C�{.@.�;�d�w��0�o��e�9r�eʌ)�W�B�K}O�7�S�]���f��C�:����o��7r�<o>o���0�`�k�l�/�����*h��Fn�����ɥ�|֖�2���of�!��%%s7��j:�sf=T��9�m��.a�.���-y{b���mND#;�'��j�?d����~���������~�(l�X5�hW�K��2��:�M}/O�ye�d�E��g���%�i��y����F~s7s��4	^�#P�5��ς Z*�� c�q^�&�pŽ:����d�I�o�6������t��.�zHzÖd����[VjW%d�-�-T��Pd}MҺ����d�Q�*�I�I��/��os>S�l��F�Ǧʷ	��/}7_ޭ���L;TOy�.�(%6��ভc;, ?J,%�N�F��h�u��L'�����c��(5���U�~r�K?�q;c�;�Iu��Nj�A"�~�H�mTT#&s�^&���E�S�0Mg�:�?ѿ��Y ���~�K��"���Ľx�4���aE��9��[C,�S��ǵ%��#|�ɀ���<e�O��t�:xw�����R��ML���T��,��H/4H�RW��'�A����8��l�A�VaJ���D��4�����Gfzw_�}�/�8�������9hn�-��ׅuYNS0�� \K"*��$�Bb:��̋KBx�܌*w��{T)�j$.�8d��[��ߍ�}%�96$$�Z3Շ�o���� r��z���~$��p��]��c�M����`"0��4����sg�1����%�p�sb��)�@��]��u�u0��nL`����iw�!�]�u9Y��m��V�#�p�	�pZ4�����Swr4�C��Y~,w���ŭ��?'Qkf�ـ�o���4���k9O��ο^ �3�����[���H�uͽB�0+��0���O���^=.\FlN��=Q��3�)D��||����Lm������>,k>}LE��ئedR���}#�yh{���Ze�U.�ɮr	�^s�r�m��c��.���8x�hR�	��8��i�!gJ���u�'�?~�U�y���y��}5&�=6��_
�ߜ��!+��4��m|�Yh@��t$��GE0����`�#{�$��t<�.�o�h�U*�I)[3�x���2~/�|&�j��Bd�vX� ~K�~�}���- =���@��۲��>n.�UW|E|J��mL����E�~hXٗ]��؜]��`�xk�������!�E�7�6���Ω
l�/��7�Nԟ�R-�I���-��W���7B�����^�%��3�w�~L�����g���䕧77a�B֥|�