XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5#0*����寣B��� �گ����r!u0�qd6l��mG���О#��;R"�XԣU�����fl�������d�-����%@���jk'y闷�����D�Z#m$�uQ�;GVI�8\�O6,q[��p��$�H*�Y2QF���[�G�e՚M��c-?�G��ǽ ��4���N�/�b^�:�O	��2��|M�׿�S��>c3��O�B9�yWɬ����-Y	�w�@���']b�7�P݇�kL�n���$)(JqG�_YW�W��;�/!)Tɞ�J��Yb�K�`E\R����f�C�9l���9pܽv�y�{�J��~zL�A�o:O-�0|6�''px�|��r~���z��ЊQ��T?�.p]n��/V�ƀ����K�1DdN��t�O7���w�݋9�O���.=�烒� �wŘ �V)�1D�;�9e� O�ﾩ<� �_���QKZ�#m�Y�7*�PXKX��x��������Jwt,�����g��N�s~	$eJ��S�")�b����*�m-���Du�r�+���c̺4?l�3����&��RO��I۝ȓ��s;���;��Fy9�0�c2�����k��@��F4���1���h3]l�q���Z��o˗��<�ۓ�?(���X@���u���}E��ud@��X"�'A(����"\d�l�4��N��RN�º��%�5�� ��ws�F!{r�� �ȣ!�$���?Z��'����ǒ_�
�j�T�s�Z"�*N��C���$�XlxVHYEB    62a7    18a0�{<!��b$�+(l����u�@(dw���[ȡǥ�w���n�.z��̗m�����a �l@���-�((����ēOL��L�b
s�f�������6*��8��I��cǟ��Wk�	�'���f1�1C���E� �q�΂)[��O��zP
����aC�2r��憮�~/�oS�gB�֐bggk�%�p�j�ȭ�'�@:�g:O~gz��"f�K	��$.s'�B7=	�z�.on��Q,��~�a��J�[�8V����,ߵL_���e_��8���X�&;�"�N�	p�[��n��A�a��9!�-^DE�����^=�j�Ao�����<���Z����N�=�S/i�g`���g�_�a�i��	&��#�9�R�|6!��Zދ��rn^Y�)|-:�bV�a�[פ��9g��G��?�f���z/ہ�O�̂K).h��e]���?�$���E���9�f�q6D��������$�mq?�]��!{����r�	Ӕ.e�P2��[ ��HZ=�~�q.��X�1�9B����W9#�j�,���_�>5��u�؀Y���>2�d3�JhQ�Ej#E��E�hK6��wb���Z���B�]��'۽7�¤��>܎њ�`��(A@��?�^�$�8<_���Q�r��T�ן04���mr��xN.�j�Æ�Z%�0\<�j���1?suGQ]u<KX�a�+���Z��T�f�.|WY��T[&�z&\��)�(7��o��3��$�5Jܗ�S��Cw��JDh=2�H�`��w��Fꎎ���k��Qu�Izƕ�����U�;�+�'ց�'~Cv ��7��v
�P ��ng�ܝ��d,��C�>�"�����S��� A��O���r�{ɽK���c��!�t��H-RQ5� x�����{#����A���0�H��A��1�UΛ�[9w0�\\�jٓh-����ltw��	A��W�i���y���Ϛ��+�^P5C\�Wr=�e�EJ�2+�?1"���G��!�O%�K�d9�SGbMG\Į�l:��T�$b����:c�	�#�;1�5'��6����#P�.<��ɪ�?��,u� �	}���A�p��M	���ڨ����;/�X2��R�}G_o��IY��3�T��]�R��7�v�(blG��R����7�/���ɤy�9HɲQ���7��-�x�1<���N�2���xG__��.��rl��H5��~���M^]��q�5��,V�ˁ�\�j��Iodw�ՙ�Z���� ��I��{�0u��AA�hh�_f�Z8J��VO�^�kj�T�qXBs��F	�W�*5N�D�IV�c�ix!�$�
�F���E4!N8�]��O*xV]�ҙV����0	]ox�;X�mjhα����qI�?
F��D����
4����È���ܣGDPF�)�A�2[��	q�M��;t(ϲ$��W,�sO�����e,�Pol ]��:�HCd�c����y�6'�}�����G�F��d[��?RL��/�Q��3��	/�A1:[�G��B��>��J��XZ�l��#�$��T���Ja!�ZMvI;e5T/R�6#P!
o�D&4~�:E�+����N\ڿ'o�q����P�)���{	�}䗪�i��<�f<֣�S6��D��uH)����qq����0�B�I��V}
kIm�9L�.~�i�p�f>3��gMHy�4K��z��&�iA�$ב;����̋�D%��`���h��;���ũǫʔ(�!���ҋ������Zs��9(�e* ���5O��z��PSpk�l��̛�6��`:�3�����U6B��l���"�X>�����maj�� ��p�s(";���4-v)�*c�L�P�O q$��Fo,; �|w��X�R��õY���h������[hI�w<�_Uv���~bT#�6�C��SĔ9�9Lg�-����s0m':U^��^���u2�Ǿ%w~eF���s����
#6B���!���v?
���l8Cr&�Y��=��ks6��~M����tn۹�:n����� �F��OI��F�g0�5 ��]���P��uvQ����o���[ �֟���L.œސ�MjA����m��Q7�2��,���*�#���H�	�%���F �Dg��h�����O�w�# �{�#70��ľM>�Ő��V��ܳ�2���}����z�4[D2���[�RJ5v�d�=H��!3>"}$ǀc��=!��*���Z+��7��];9��ҭ��d���0g���ŉ�~�΋����4Լ��8�t���W�ܓ�V��m��濈�z-_�:K��/2<�`�O}��O
/��������J�Q$4�Ұ$�Uٲnĭh?�f��z��Q�N��{�\c��l�ѿ�#Yw�񒇻',`{�]�� ����|��Y����	�@��Np�E(���u�j�ą{�2'À�U笆�b�1q���y�B�J[�)�jE
�j������ga�<I*�F�¸�c����[�|��Y�E^��<#Cn%�����Tw
��k�Qf�ZL��W�C���ٜ��� ��S�?�:���}�أ�1�f�˺�,ݻ�o�w��1�Lw��ѹ�wL�,�QpdѦ�����/!�����39fP��-4D�ށ��ٹ����7
G"JN�B��R�A����K.��V�D�N������O�;��q����[��5���c���IW���x+W�1�!��XIu�^p�Ko4��g�������7nۛ�����u�Ԏ�&�s
�3� gks��ʫ��K�o���6n�y��U� q�|����_*���sꐈ9��O�/�9���Y��s����M #�8��ΐް�}���4,��7̕�!��4J��\kERllɷxN�T��Ҿ�|]fKX�L���)��ѯ8�*!X��_�-*,�j��zg��x�ę_8.bQ��\&MZq"���7�n�X�2�� �~��G�Tp%���&9CH=Ѷ��� �*֞U68��C3����sz�L���+��0x����Km�I�h�ٺ+��̱`��� !���!�e8[��{?����ވD��;��61�A�q�f���1'��"C~�����\e�Gl��{�y��z-��#�I*phA:��`��4����[�HZ�Ҫ)!�dc$�*p�O��	 x�_�7�®�M��x�ST�3҅���H^g)'����o���3��jo��ޚ�������yͻa�6�P����<��x%cx�����L����-���pv������c��\pl>�)-�hH�o��j��:Q@�7a����8����Q�,�+��BH~0z���$�ǔ�c���qO�{d�x�&�r���d�y��O�����|cl�,�i6c��Z�C��M��p�j��Z��Sɉk�$�8�i'�ca,�5�e]+����7Eyk{�G�?]a�����Єx��?l� ,F���oU����ի֜[(��R�U��������n�3n��*��)I�D���^�;��Xn�	�,�}�>sP)��Dmgt�ﯾ�g/�)��"�ҧQ�Uh�d���:�u�����֯��B�|c�WL�Ƨ�{q/��Z�s���Hn&�^Pw����Qǭ�m�+�IF&I�p�ׁ��o��,U��ؚ��mA�F���n1�$6��������с�����`1Q*'��̚S(J@gX�7��\-'�j��q!����I��M|�|�C��~�7T�a�R0�f˯B3K�`�n�O%B�z�r<�8L�Nᓁ�j�������Ia��#d����I9d�����0��|�2GH,���ND�M�`b'"�n�r県κ��vFv�\tx+��`"��o�EՊ}E|�Uv[�b���~��.�o���l!�w�VN��Z�J�-#�ҏ01�#�L�����2c[n�5�
�����*s����N�U�4ү��x�:L��u����[u`�?����:������G\�lC/�=�)BL�1QA�����t�ez)��u�X����7��Ϳdl�W�o�0�6�)�J��3v�ܓ���uLXRXb�",;��Dhg��c|���ti�H^kL������G�B��*e��6�iT�����Go6��	o�k��}�:�v����G�Z���侹��|Þ�G��x���&])�\�v���e���G�}:�L��Q%qG�=�8�]$�6��QÈK�>��/@%2�K�}K��7):��������ӭ�;�2�"����t4�*�AM>N4�9�ܿ��)����E�a�:D1�c!R��c�n1E�Ǫ�x�=�A�c�5���4=��a�������Ki���Y[T(_⃾�
�jG��D�$�i��k���f��"7hJ��i`:W	��Z�-y<���=�,���'�����c���؛zЪ�Gon��ٔ��X�>{l\�'�*(mc�+M�G��t`RF#0lǱ�-��@�Q\J<�)�],��f#�#�ee8<��'w���E��?��>��t_$�E�G� �]/��VRt\��O�7򡐐*�r���4,�>�[Iտ
��M�U�j�W'&��l��1��~O�֊cF?p̠�U��(	�O��,Y���s*�doo���k����b�����{�_;��0�I+��0�͉�S@2o����W�'UQ`������'�&�4
B�}*C��:|���RC��'���?���eh͒L�]H=R��;@�Xl ��p�����Ɉ9��0ހD`��a�2|}���x=��2���N��|5�mAv�v$#F���cel�	��٘b�
��z�S:�B��#�k�|�;�nh��n��M�e͹7n��,Lڀ��ƭ 
�%� _��@��V�����㦛}Jq��-}�(�_ݡ �С���l2��2�-d|�LRg��<�j_���BEr�+ȑpK���9ETLDb�:$�=گ��r\���h/ee�7�e���M$�>��.��1"%D��^��݊�B�ſ�
w�:�'%��I?���M}".pj�������yQXF�Ϛr����K�H#���bB[�E���8�̯Ը���+	i)�m�m�5���bu�\�h���L�9��=�n���� ��{������Q�rH�9�� [>��`���^�{��_iU|r�T�d��<XK���*`G����m<pWd�0��+��������$<����5���"O����r����7+�ߪUΩw����F,����XH*?Q6��Vy����&� �4ֿ�/\�6���%I#7���	?�,��r�:3a�(�i��J��j(E�j�8J�'ER|�c�s[)'-{���J֍_̕�u����H�e��Z��!���P9􇈔��c��:�?r�p�����+�ݲ���L�@׺�'�Nj�Z���y��u�S(�+1p,��Q�/�*�{y���I�E�������4���DPE�x)?"��j�T����%�9^�	i�AG0���%�N��*hZ��|�(�i-L,������s�*c<�!ۑ��n���>�|`5,�\vga��2��i#aoN�^CU�sbGrE�=�2
ο�)���Y������EN���_0�:z�&jе���1�/� %g�G�ddT͆T���O�ȆuH��"�&m8c��a��A���Zb���DD2�K*�'Cf����D�W��]�1��������C�:���S�<�Ƥ�	��GC8����yP��qɕ�q�l¦UL�dt�W���;��G�0�� �m$4�j)�xh?;;�I�>�@U�w�	�?=�0��me�j�3�Ns�Zv�űӝ.�Wx`�;���+��V�w���1��p����d�8�k ��� ���Fk[�μ4<��pqw����2��_%��]>�;���?@���b'�*�-�B��+�f&���P�ۦQy��J�xnDoj=��YBwg��`y��3"�i�����s�$��n���嵹ނ��
��� ��b����%���h�I+QX�C�hϡl��'#0�G95�� �N�kb_}U��֕z�.)ֱ����F�L�;��M2d�igpe�)+P�����{��0��e�m$�z4k��@q�x$iJq�I�����:�N_>5<���w�}V�r`C�^#�Ð�ɫB=