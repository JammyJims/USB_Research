XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	�"文%��t')��K^�s��0\��{�:L3c���[j���,��1F�醙��4$C���evޢ�y{�3s=�����D�ҝ���ACn �d���`Rr�o��3�S��M�a�a�����e2����Ja��AF	ռ�ѐ�:@h�,�>�l�B�b-���9W߂p�16:+��]��Т��4n3���<@���6g��5���4o����,�/<<�C,f}���|7��͜{��,��,�k������v\I� 	�8~�E�=�W��J�����8�m$Hj`*zU@B0�ၪ:���E��Y��ū����}�p��p_�Z��T����Ӭ3��L1��u+Ps��5�]�5��yH9
���w�B��n/C�xD}v�s�Bp��\k�������!�d:F�L�)�$It@�f%�n*��|R�Q4*��Z��c�A�o8�-b%s&Χa��3�Ӛ��F/���%�;aD��t�9�D�Mc:��A�ł	�se�KNLe�5fL����UR�Ύ'J�H����}��3m��A�Q��k��W�l�	�k�(�A�N�B��L����d^6����a�u1C-t�~����l�j�W~A�L�`��(��&F�w�i�A�-�Od;�� <��K�'ѴIk���x��tа�qh��d��?���fl@i��lX~c9���H|�GE�?����s��🈜�D�Zyɳ�W.A����t�7�����3]h}2�������iC�I�XlxVHYEB    5923    15a0c�t�/4ƚ�a$�>��S�F���4+���ܽ<v��{0Fm���˜�c�<�[�������>û���Rzx���%UM��)�X�[��5:a�>;��_�(��3�s|p�Ld�{T������G1aR�T��Rٜl��a�=i(�gMmC��G����*[�m�Ʉ �|^�<h�� ����qMſ!�浰5�^��l|���5����^��݄|
ӂ̈�ŷ�v�Pka61�]w�W-n�?�$ݯ��5)ߡ��2��tĄ����V GO��;%��ʭ�f./`N5�� ~[�����9�F/�
�i R+ٝ[��x���1��&�Ũנ� E��`��(>d8S�Q�S3���� ��T�����)��)�	u2�C4\��d�gX:���ц��
�|/u��V/b!-�)��/�D�ӗna&�yP�;�u�AX(���d�baM�v�9�W��J�2[i��*��e���v���%e�q���e��I��#���M�����p��P�9��-�ݴ�ĐO����-��h�"R����qG�^�3$;k�I�Y�X�_�XLz����%����(�_�	_�>'\j����3�e��{<[�R�`�&%���(����w�%M[����{��J���o#�/S��Q���$�{O�{w)DZy�KFă"� xe� _%���׻�j[�$���oy"��)�Y!���9"dkPp$M��ו X�@-��؉�~<ia����a��kx����k�3��A ���<���،���L� ��Qp]uURZ���Go#'g���D�"7,��P�BB�<�H�kM]��9؈Z�0!3h�o�ͧ�alM�`���A�g���P��~�$:�a�(�Z,.�8��`�So��/�5�ʴR���e�`����Q��B��B1��f24�@��q�4�Osa��������In������ۥH���'���3Kh��nQ5=�d��[�j$K�2�<��'���RZ��zⰇ5��o� Q !w�xdw;5�'x��6�[��PQB�z���;�`�J���!�{�F�/� {�����T��I��
oɫ���,�"��J'���Ees�]�$fw϶��+�2���<AuB�a.�a�_sM����8p�2�([	wC ���|~4|��{���˅C�|�����i}-����Y̥(R8��~�A,a����>���6o!&����ɲ7�0,藺"�<W����W��r6��f?�bdL�ppqj�ρ�����tܰ�x=%7�e4�a)���q���&]�� {j�1��� v�!h��_�ܸ�/��b�%$�Ss�kV1:qW��K(��C���㔲�]��7�$������{�AE�WtqU�;��򶼹j	T�Y�7l�oJ��.�p��`K��ݭ���|�"pt�Cf���*;�V9��:�bo�d���D���M]

��#��j�)�?<�f���z�ek��|��`�}V�L=�}i�B�����d��s
C����L��'9� f��O�?��\���_�+�t�O�]g
���{0r�5�WU1�&V�i��<��.�r�a�d�k1f�{6�s7�@ӹ�F&zf�Sjh���hr!�����%p���hI�:҆|-�vw�d/�X|���� ~4
L�}��C����|v��qt���$L
��<[�^����&Q�K5r��q�H �=��(B"D��3����=`<��S����d�/��^Oh19�]�2��jPzL0�P��h�Bz�_�5fG���딿��:ٟ2�0L�ܖ�7$�����EH<Gax��@���e6�v��gG�Z��cz7͓�	���M�~��E�C�1.�}�B�逶h�n���9��0o3�,F���QHթ:;�����F:ǸF �y@��J��g�0<��CS���נB0u�=�Vb�̤�:���{ao��e���jH���#���S�+���٨H?$BqG�F�Q.��<�����f���C��m�|GD���[���|d��K"��E�^li��
A�̷]��?��ش! ��� R��֔�ݩUr��]��L#y�J^����wFڣA��%X����{f�A�;V�켙����� ���z�կ� �oc�2��jO/�(Z�4&����%x�c�`&����������e&��^�q���`1|�=��kH�����a��Qo~̍o����O�}���w�h�V��l�q{Əv~�x䌞SY�7�����w�lk�kR�ӆg�a����}�W�_�ȵ��`�ĝ�e��}(Q���ӹ_���o��hȿ�c�GS���o��x���)�B���XU����N����"�f����]��p%�D%&_�
ǟ§��>� �9���*K}K�H�>˙u,N�9�:���s`�ʆ��ڭ�=�W�J1m7�-K�Ɋ}���;���
�g�k:��rֆ;T�lw���Ό�����I�nY;T��I��J�r���c��&p$�	_��;(���P������cX�����8��h*m�3����׿���:#j5Hy�.bT�v<�
p���w���2���Hs�x�z��N���:H�¦�C����m���_R�[;a�7e��$����8ԗr!��ě�7��"���x�w<��@"�}�A��ڢ��?>��b5\.	�?�T5i�a��"���wKѼ�a�3,�d���o���U�e�M�y�� ���S4���X�	|Xnemo>'R�0j9�tu��~��M��0t��	��ti��hQՐw곆�&���K��C�y=Ō�?��vӗ��u�Jo�"C����%?�T�y����/��$1!�>W��#�*S���Dܬ͡V�����i��Iu���Hl�kY���ֽ�fJ����ۉ�dn�(�@.��P��u�]�{��b/�ǂ��@_�T��0�T��t��L�ɡ�ѴbP���Ң���a1�"����XD�js2[���qU�����9��Gđn�.F?��Dv�?��2�^��2�uA��qS���G|01�@K�;���D/�����>(`�KI��ݒ�Ɗ�.��D(]�:(�O&T3=�o������������G�GP�4y�4!��SѼ*��:�8f�JN<����~L;�;����q�ƚ�����z���.�s��O�h;�3Lث��v���㹑Zx���N0u���d�0"P��WOY�m��!zV�N
���?r̅��,�OhW�5�����b�]/%R�=o�v�~by�®�W�hp�u@1��_�5!�`�gWɅ�r��ʍ��k>�RTC���c@$G-�����j)�SyI8�ƕ��},�������RR�0���;�da��uTG�xN��xON=��e]̞�I���	�� ����[z�3a���F�~���#�[�8a�vy P��^!U�7ǎ\1q^�	���̨dp�N�f1(!=QN��u��j���!���4��Bv�b{+h�`�Z_��������ﴳm�N�l"Aī�f#9�H���d����� s�x�jL��l�3�
5���I^m]惴��>�#�q�%�L��l���u�C{��ʹ�Npy
W�P�?5|�E��|u����N�w���ُ��<BC�ب��{�"g�簣��E��q��xU�����z�Z1�[~�ZuV�n��F�Zw������K����|���T�E�}�g�yA�^r��ɹN��'�;L�ߒ��}�'A���)%P#YnC��B�-��y���v�"��3��*�h>T�>$�l��2(MH���������T��6|�o��k}�܂eK�ZCE���
�e^�+}���cpv�(/��!��Exl��m��*;�n��T�\AZ9�=��eG9�ܫݽ�n�By����aw?��3�)��<$��F>Y��cg����nF��V#u�HLSD��t�ר��4l?f��g�Z�V\�\1t��wN�}��[5�0��<k.[�)gªm�&���`כ<��������!�����`��B����S&v�0�Nc��js�^J�*o�ԟL�B��$�jc��J�WKӁ�x�h��2�$"_��Ab�|��倩<�ɥ���a:҈��7|����G�h�Σ�O`������mr�5ӑMWåŪ����t����!�V+- ��=W��tW�ֈJ�7��W�Y���<T������H�*�/I��햕�*!��Z�̥�}'�=Q?r~���H D�_��
(��!Lg����i ��U�f��>ZF�MRg��m�&k'��|��=�6yT�{s��~m������$�i��U���z=��oG�o�7��g�ܺ���S (G�C���^�)�a,?��u�����2�!�BIj��<�*��r�|��愪��bF���$�X�e��"f�`�듥��N�pz�Q�\r
6*Ԗ
thph�}��3Z��B���9����>hZ�v��xE=E%N3��o	���p1_�8�$'�tἝ�R��>�Y��(��K����>����"qS1���5��Bn��"��r��UY����������;qu<v9M�v�.���ޘW���i�� eKJs�\yQ��U��r<�9���R}I�����.��
h@gp��(jev�q�Zz�[ M���u���qk�aq�I~�j剼<�Fe�]�,�sEᒍ����L�����Iaj�o�K�;g��~��?W*K�`�kp;�� �`���q><���.��Z�)�WQ,���~c_�kK��Ij�P�6��F��`~��Qk��sld��j��g	_��+B'�WJ��O��'[�U{�,��5cBsS�;��7!����A�8NK�����>j�Ђ��*ޛ�ٞP��ޏ\Q�(�Њ��*⼣,3p�Q���D0|I}���f�KR�� GT+��`3a����z�1�ߎRޭ��W������3�,%\
YU'�NO�8.a��a �A
��<Z�R)c��͡f��I��V����ܲ�@���!H��j6��;�(!�-������T������y>w��ɯ���H�����J�J���M���+�����<8�8`s�w�oS��E�&�N����]O�ܠ��:���&T��$�Q�OIJa��è�	�w�jCZռ��_�2����}�VRXB�=)^A���;C�10Qㆮ�R�aX���W�A�"Dr���w6���k�khL��Vd��;k{�s��}6X
���$�][���͇L��:��h��liR�Ji�V4���y��fz�Q%�
�ڄ̨U	A|�ӳD��:�O%�|��Я_���%�N�N��D��O�ʆƷ�U��b0�N�W�3����΂ci�97;w^�T͋���>���@����9�e0�.:ʒKvFĔ������J�5-���