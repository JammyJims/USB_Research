XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���3��Y0.�c��&��$-����֏�6*h-���z���J+�WҸ��~3�_P�5������8H�%���7�z��)D�c�u-��� ���Sȿ!�0�0^���;�8,���X5�&r��6��ع�?RJN��&
c�4��w�_|6�,�;�|6�M� q1l�-y[��̝G��e.X_�J��`�B�6B�X%�/�G�z˭�K�m,�HoۿSeH]e����n!�,�ͬ���s{� �9�F}G���o$5������g���wE_��CO}�,�
n�(@*�3�ނ+B�����rWM|��.�[o��'��
T.��Q\Dw|'r�]n�bjV��{�ށ�\�������❢�ێ촮F�0��8:Ξ�1��
eY��w�_6u������y�;gE�8��++���(eDi���ԪUZE�%���U�w�٣dQ���?�Wjީ*��� �2��I @��WAY�J�~����������}BRdG�?eQ�z��G�Tațr6�оK���iT��5��a�zA|/}�L���֗ƠQ�4\�4vm곿��5����;���L�4�CD���ˣ،P%w��	m��C#�
A��L���c��Kk���nG�*Fx���2�b��A
���%^ά�{���#$^�d������*�D�u��,l���+Y3�f�9��)L7k����I�@&��!�p���]�*79��YJ&1�4�d�hm�]������l�h_(�|�X�����PYXlxVHYEB    59d0     b80��&�Br��,�-���,`=0�3���[��N�υH�y\��g+I�pt�v-�޻|�nF���ZoJ�m��	�/�����T�E���ܚ�S���2C���
OTX�Jʨ���\�u�8��Tn}J	aHj����[����c��x��@�B��Y^����O6��jD�F��˩�<��J&�.qӜw���ō# w�Q�vd��y�[ S��]�����D�F'"��1J��?]��S��2
��[uxz_Q���܋�n�|#���-V*��������ٌ�#������S�fG��-U��~�����YsS�_:����&��Rȯ&3)2�PM�:�8�3X��;�~��R�<�ۍh���>
 ��^h�X�c�
���
��m9�Si����Y��Up��aH!�~b_���40	���R�?ϴ
?�l+<~a�J�Q��ލ�.�铗�G�gj��P��5�]�W.�����{�*�uإ&�;5������L�HK~/�b�g���LP�+D��;�V�&ЖH��v�P���--��"�ʁ M��.EK�m������rD"{�.bd��lp��;�;�$���=��"�]���(���~������M^8�Y�\�$� g���C�L������q4�q8���Y�MM�9�����M�����@Kk$`����{I�BS���%�+D���í��؄)G��]��W���ŅW:�G=Uɴ�� P�"���\��Q��������������)gw��$jq)~��{�2���ϴAQԒ�0�^�E��_m6�
�w�a���-��v�eG�D��gk�8�/x�;
�D:i�n�x�*��9F����q��G�4��&"�1}�4V��u
��r]�h�uaT���Fm�����Z�]G:��V{d�����a���nF��)3�݀����=0%k��EN=+L��:6+���}uF=���uf�&.�d�j��ِQ�5��o���j�Y);Kn����c@#��|9���JI_;.	��eW�]�k��u�վ�}Mea[�DMP��HaԥQ�NR��jb}��BaP�]�LU �� �\�nhy������u{W1�1S��T��1����,��>S���
�����%Y�\H�+B�a�0"�Y��RB�G��Wl"[�%��5[Ǔ��[��]����s�5�b妻�<>�/�>"mG�XX9n�v����q�u+�D�\�^��6��Ia�h"IY!E��HGk�z{���+4Y�
Ye�_Zt	oVj����iQGo����<�	��n=�P�Q�ǧ�^Ѷ}E���*����^(�d�BQ�:I!�4�.��((9"0�d�7C��������s�����h�Կ��|�����k�A:'X�\�2B +y�pİ�����������N�a'Kjl�3�V��v�f=�kd`�N��zT�ϑ��<k���p�_����Ǐ��Нٰ��b��A�8���X��y�<��DAv��G�ޤi��/$�Lק_���$�qn�l����E���7���w'��$R"��>�hX���L��i(c�L�ҹ��ݧ�w[�RwO���!h/q�b���p�~UM3	U��#���������|$;�Z��XJE�^�<���`SI����h����8���=����(8r����/�ޗ����;+�R%d�"�Jª�W����gH�=�1@�.-�,8ff<�3^#�l{��	��69d�pgf�=ѻđ*V��*W�4�(��Kw'�%��A��]x��;���Hy�O9刹�x�5k���<,��sΪ��"���G�Ѯnu<�$�����vzXI�Ǹ��L#e��U�<�u,�*{�`�ʝ���k6Վ$�}����
�y�=K!�b-�h��zŻգ���FȂ�)hF���~���Dr�Y~_nd���5�M���A�������"��7�Zʀ0:�e�ר����lo*�;釚6) &׽�5��mz}�O�1(RQ]�"`��g3��$���:�ӳi�e���鿊���We{d}+T� #��P�j�ԍ.������fem��SD��qÐW3�K�/`�E��Y��LݩFb���>�&�oO:"EY�JfeKix(*���:�]�yk� 4��o����D����������,<��}v�Ȋ	�c���Ix�x)�J��҇i���&0�~)}p������֚���S�;.��J����b�oJ@qbU*�L~�,[�\@P��臁�X��!��%�5ժ2͘P�(ǜ4A�:��/����s�#I�aL��~�U�T��qƉ��q�F��^/��g�4^K<k]UAf����������	 �Q9rzd�	�O&��3���۸'L ��H�I��d%�_3�M^{T��1�z7L��㊠������Pڤ9�sF
�%Yk��*��yg�[���� )�v>�$��#��."�v� �D���d ������֍����x�N�����������x}Mef �:�p�YVF�={'�_;�B�c�A:�`�Y��´㋻տ�J��j`(�?��}���1���J� �C���>s�����8`����_}H��`�$��,����.+�N�3���yY�jA2H7pU�8����4�1�t�c7D$�9@��$k����s3�E5�D�|����nh��8�bJ�A!����S�K�6qcw��v���u�7?��!m8RRG�X��ʚ�5�$��]U`���?� c?�ǵV�E�k�S�����b^�Kzd�d�_1��3j�g-#rك��{�\����w�J{���
�,���E��}l�D�ŷ$j���GQF;OH�i�Ҡ���/�M��<J�r��x�����wלq�i@����9��_V�{�N��Pz�