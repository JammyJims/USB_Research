XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���?��Ϭ�t��jP�ɇvˢ�C�-b�����u�g[��l�*ɸ��U�%��`����\�3F�i8�����©��{��De�28�N
)o���f��ĝN&T恖�Xt��I������{�=�2f=��\�k���%�i���yh�Q��Q�_���PT���$,�
�K�_TXw��b��-�ó��B��{�M����F
nR9f��A�E�Y���8�Cu��]�w�H�(���{������1���F��ojԑ�MYl�/d��r
Y���(�K�Z�����j�-B4Y(��C��L�;;<���<s���&��n�U�~����"\Q8�h��\��:�F!9_�� �j�2K���㚆�_��²�>!}� +�лZK�g��Vi�R@1���{^1����炦2����	���J���0���ƪ�*�G{c�%r��f�4�b��S��l"~�*�����t�݊PoV��+p: XӒ��	��U�;E�t�C��~Q��pᖊ�F��dl���/�@DM%h���uO�:�H�{܋!.�h ���w�4��ww�\�Qo�`˚��^}9� �J9C�R�a"�\l �|/__f�*ô��g֍W&ۗ[�P����>op+2^�J�W�[�S!m�Vc�����C2�<�@�k�r�'M�zMHF���'�T������Mf'��_��T��Dp�?�z����J�������ɦ\zԛ��y++���$�WZ+y[�ĩ�)�I�!�H�B�XlxVHYEB    9981    1f0066��( Ő3��� (n��gl'oc%�u�i�8�?5u{�e��Z�#���Ф�
�Wf�.�$�=8���]j�,t�a��r��o��93lȎ�Gf��3;]��z��;'����`�Z���z=]};+��I5�r�}I�H�;�܂���ʣI�rCڣ�P���ֻ��`��I�D5Q>��ި�ÃL�h�l�m�=o:#�A+y;yE4/�0a$�
[8>ѵ��=�o��
�]8U"�ܘ��O���^?����Q�ܕ � G�0Ϟ�`f��~���,�I��c��*c����mϫɈ���Ϊf�cT9(�/�|�G�r�Tǉ����W���.��^r	���H�}sK�v��ؖf�]�j�ǈp����"��{���t���GM#�N�2�ޟ�4^f�#���"�~!���} �u=ͻ�Ba�B��=F�:�7 ��B{�lmb;�g��|���0��EK�kY�M��0��t����T�>t�T���UW�4m�51�٪�x���:ʂhC�q��!0��,���ֽg���ǇUh̀RE<������N(T���&E�e��I�|E�_=�����Z��](,/+�콠Oi�%XN�V�����/
w��6.�<�nV����(.��"�e�vV�X��n��,��]���$x!w�8��5��PJ��R�9U�m�A�r�a5�P�`��43Y�������U#�n�M�(���/��J
SV��L˙��L~h�Mˋ��J���v3�6`��kY`��y����e���Y5w~��~�yf;�����!ȳ�Fc��a�U*oƔWaMWȖ1�L�P(����@�8��9�"��1|E�O�2v��y�G���~�#Q��h�u/|;����cX�!��Di�Q�gV+K�2�v�x*�G!CO��p�����z���U�]Z~��Z�����Dtb�Fr0 ��_��ya�Å඘q_�b�k�9v��dC���j�2̕N��// '<��C���&zp��>���KZi°��u���R>��m��<�*1�aH�
�`�����e�03�Cfڴ�ꬆ�Rrw�D5�Ӭ�v���U�X�^�j�����/�f�r;�(Θ�aGK�q�|�9n̝y�#"Ӆ)(%~N��'�l�v/�����}�|���h�,A�pE�Ǡ�9��"��J-�"�o3f����e����?j���_�m/J��Y���.�n������R��B��h�ǭ[G����Wu;>dH���'���f����Y�؀F���ە{����Ad�K�造>Y�3���9w	�B��>�(Zrr{�]yW��|��!��gǥm���f*�>���I�z�@�rJ������(GS=�Wg���@9*�7���UF��閵a+2W���y��h/�!�*��s���C��V�����η�*�H^��t$��w�׈�6?k�Y��&�Չ�y� ����Ŭ����v��lz��\Mk$ʿ���=eS�9^\��#����B">���䌙�,�WF���km4y<�;XӶ1Tْ�E(��t�{yI�i�A��!qè^<��i!�[ԁ�.RB���M@O�*`���6�?��bt`w�>T��3z�x3��S��J�}>�*��U��^�G?g�q4$d��h��J�AGGPw�e��T������h�W\x :�߮	�8g�5�;L��~�r9���'��Q��↶���"�d_�p_x P��J���G�An<�Dsb�6S�]8��p�M�n?���a*�^�Q�亙Qm��"'5'�"'��w2<��5=��G]1`��@�6��UV@������k�h�� ����޳���.p�<:�	2�W|�\�9j0V������0r�RAtN�����]K�H��J(�x,FGI����
\�����z��"�ٮ��v��!n`Ӱg�KI���:-��վD��)3��8���l��w��l����Ӵ�ހ��W�����o�&8��#�Z�ʬ����\݌�?�/��K�����]�Ԍ�󧰒M�Z�$���=$^H�v��w%���K୎k@�C�l��`,esP.�Ԉ=>�,v��t������Ѳ�gD���^�͑,3C��dE�٭O�����Ek3�\�"�o��u�2 c����J�%_��{Y�Kk/�_�#=���%�F��ȹʸ��jfk�f;ix7�s�rI�@1L+�mή%��S��M�?��X{��{J�'!f}�.�y����5 ���� -_f�D=H�eH��lWHx94;��۟�=|�r��s�6`��"��/��I/RC���w���j�Ȅݳ5Z�ˋ+C�-k����oW6�Q�@��^��Y����_xq��dY�w��$2���).�=J�ϸ	��~���*)3�d���P�	���t� �0p>��l�g��6Q����vbEj,n\��%9�%��Fm���ء�=�z�)
����_S�k����2�}�-�;���y�����D��Vv�z4}�9(��^���2�V���K��:��L-g6Nn�.'�������X��,$0c��≺iE ug�7�~���@N�nz/;L��͘�����⿏.��erb�t0BW�5�Կ�&��O@3�zs�CcE������Qoj'.g�
\K�yp[�n�ެ�{Wwh�����+e8X��ɱ���6�>��r�� u@^����sV��/p���JX�<פq$v�L�����9d�'�69͟�����dg������X��R�瓽�~�4�$�X�����'-�
1�<�U����o� |�e�v�&]	�e�~Sܰ����鱬���X�qOkM:��#8�=��Hn��&q(|�1W��{,l៏8��d���^?�����$O�m�ؙX4i��6X�8�8�F뎒_���f�CN��ޕ��Q�Q`�������o��x�/���[��_`��D��j���^9���n�S�Eͻ�N�Ӛ$(�$F7V�Z�հf�<�.�_U�S��q<^=˦m>_~���{o����	��嚙����;��{��pr��z�s�xD�n��O3RjK0���*%� ވ}Rh!�1F}�3�K��q�����^���ą"l5!
Z$�߽��R��9�!�i,�qkG��^Q�<_iR^��J��`G2�=v[z9�AS��"
�҅,2�=�S��鹩 �f�0�$���ܪB�|'R�^�o?"~ZB駣�<'�*��XP��AH�m�ɷx���e���n�]�S�q(Ed�j���9k!�U��D�m��r�_hF��ҿv���5`s���7�`���v>أ�|�}t~2	V���o�:��F�=�ˠ$?��e009�G��q��}4<W��.�{Z�_�3Z!�D#o!�e+i�ڴ*&d,Z	��5a� *�=y��`V��:w��|5*ˋ.�7��{C��?\�=F������Hn�h
��]:G%.�&�
�g*dV9��}�M�pB�w͋�����R�Mj������Eaۀ(�%9�%���� �ˢ�(��%t���c?LPL>e\+W�3��'z���� P��������#�w0�rz�d�ԔU%�#��)T7Ǣ(,�c�V9Iҍ��%��i�A��_�q�w�m��W�d���z�8S��2^!�,���2�-ֆ�1���Rr�x���:"ʴ+�dM&L|wy�dܯ�/�zh��,i���~��+��_���:Y�la�qp��ϲ��X1Ňjzj�� ���ͭ��I���m�_r���/�:�x�@M~8�F�5�=$��ϛ��������dJ;e�lPH.��S��Ds�.ednI�:$c�Eƹ�2����,c��R�t|YU/l}Q#E gJ����䧲e�p�Ѩ.��8.5b_�G��(��DM�֧D��ksq`�hz�h^�.<�j;�C����f�|���E�y`�/�g�9�x}��GЕ�\O�TRF6��+�5Gl�?��a�|v��̀b��g����v�z?��&�B�n�g���@m�8��9�)�R�  �!�M�P6�ꩶb��Í��x6,���iG�5c��݇�k/eG[�'2c��BL��w����Sv�	Kj�7t����oL��V��+�z�"ږה=�5��/ ����B��Yv ����PU��-ku��'O
�l��x��Kc���'Xˣ�E�;K��.ƕEYOD�i����yK�n}֏�ҍ��2(��\o�1��L.���geQ�"ی�q�9���;�Я��jJY�<@�D��\Ze���u����o�J@��1?9�)�.���V�-�����P�u���g�	g~���F�nj
�ܝ�)�j/����3eZy��hj�3t#Nm����D΢�E*2T@�� �)*N0�_�ht��<�
t
{�RD��r
�f��t�r�@.˰F�m���ۈc{_�䓳؆z��]�X�L><]{D�Ms�p��̒j��vS=�]7ge3�MBV�m��B��@���p����p`#tNr[f�6����8&��Uȸ!�ճGv����ym��`<��f$��/��c�P{Kf�VϧN�O�է�\!���J����Fc`\)n�6����x�bL���ѓ|h�'�j�4:�����Nr ,vn\�f�H�z�Q}*2�2fߖ���yʼF��$$j�]77��g��6�n h�Ce\7��\�T1�J������i�vbF���T*\2�=x:5��ۯ!���E�B�@l�Uk�D�&�ݚ]��� ���D�wи&�[�������.��zw���p���к#� �O&���|�s4yZ�ĸ�8C�?���?���1B��F�&�Go�[�`��������qq~&~��+��4�{mHOl�Yq0I�X���p�ZEa�[H�{�@=�HwFJ��*���'�+��Ɗ��K.��[�5�uz�7�f��
�9D�+[A �s��H^�5;��p@[o�ހZ�,ZC���"`���#3P � ؅��*�^oC��Ñ-��౤�?�{��^��ua�>w}�k�|���4z�$�{�lXe�.����<[Hs$7$o��D@�}0�ƺm�ۉ<mpO�#\��0�-L�M8"�g�'�k	O�ޏ����d����e����=���Q�(��B@�����,��ڶ�\{`Y�i�
�=b[B�s֡n��>�C-�{LD��󝌢�� rW��w;���>,��n�kA��1�c9�c��BC�&D���2�%��)~�ݸ&��[7���\�0NQk�F���L�˽�@�F-�x�`io�һ���ip�~Ws��*ZcTۃ~%�&s�qf[�s䂦:��'Z�~b-S��穬^�P�9���ֿ8�>n�TBOnR�P�#�*���^J7я�p������S2X� b���N�l�)삅��-eB>`����4 ��e�~L[�v�x�t�T�� w�:9��6Pa&�"�����&V��N���B�2�}{�<���BH���\O�(�^P$1�#�s9�s�С�(���t��ܖRD�4	�Hqm��w숒�5Q���MG���%�&����P\7x�Ni&��&8�V¦ŵ .���h���6�?��cGY�A��:�rM�M�{~58���d�;�(R ���a�-�5��t�|;�/V�[�EG����y�^��_���L�#�R"�j��bN�Ȗ���v�J�0
n����O�vz�N��p��k.�F�>�(x?C�ك�s���L��Zo����)�z���F v�@�}����μ��ŎT0�m������ˍU�zK�8�qw���7o���J*��~��b���C��-��䶌CޣD�N��O3c8u�5���_xU|w3�xRc雈&���+�+]�a�$` �3i��		iڪ�>u���&�#jjAb*>Z�M�y��)B'�_^�ܻ�9U\��T���rcE�s����.�_�0cT>��S�縣Sxr;,r�v-�Et���!o@�5F]��X�vv���I��rm�6����8Or�-�|T'x`�_����w�L/@&�$��?�S\�{�(f�Q��( �ax�;��d8�]���_�6�	�$��a����;@?�L��M�=�j�A��LqG�8����#6;Pʸ~��Q+p�#�ţ�`�T���9���V���S2 �b9Y֋.	�4j�Z���_��쿂�=��k��nx M��h^�#����]x/��
	�2�e������b�"=�6�����KMo4;�7t���x��MP��^;��d5��1��Q҂)�"��@w��\�/�y�,��DZ��2r���v�;�b�Y�� �aM�X�i�z65�n�W,`̪�gh#�Y�E%�v�,'��1�%�]�L=8L(�8���"�E�73�:=����z߰[�I�p麄Ʊͨ��N\�c�d�� JYzk���z�Є�<��ĳ��7Ͳ"��	��]�i~�����*���aMЦ��n
���z�K@{�N�����	9���tZ���壨'�B�c��2�b�2N5���đUJ����O �U��33_��+;p[ ������,HB~2���W썝��r�W8���Sє�=���q38�1De`5��ϽL�K�F([�q�e���,�ܸ��d�B����G���v���+� -���͎E. +�n������S
rK�R��8��|�0�j�
Tȭ��E�;|�x!{����mU�0���+��vz�
��"�n^.�U��1a/xq�H��$�6�<A�`�M�w�v�׭��:���O���B��� ��nح�e}�̖+\�q�]G��XE��jG|l0w��nk �.��4R_.f&	�T����	"�1F�5P�E��NSJ2#�� a^�)��`t	�^�:
��Vi�[pO�-�pjQ�beҏ}w��-&�vC�4P.:K������a���W�<��ҹk�S���πw�B?L��pt�Nh���4���67Q5lm`�p����	�ǵ_=d���0�oA�0��-%�TW�[<�tW��*R���7�,�6�K�Ɔ�;�p�V��~������5=َ�<��F�Q�f�g,B<�\Y� Q0��65��ǢKB(�Ӈ�Ghs���:7�12�i��W���S̑LP��gН���4�x96m���l�j�n�'�$7�Z���K})��9-� �9���|d!ћu�گ�Z잳_�1�M�E����2z�
�vW"]U��>��ܩ�ڿ\�����2�����wP,Tr�Ux�U�o<]����4^�!Bx��Nh\D! �!��?��J
�@�C�d��%8wKYc_��`��j2�y�"��W;,��ymf̱ co�0��eQ �p���x��D�]��3��x!l�I�QNu �VV֘Z�X�$u���Ŵleۍ�X
qJ���pjXHj�i_[q����$�:I�E?�W����W����E!�Y<���yfv�a�Q�s��f���j����M��e����;ZϜ�i�CH3�ٍ�A�\O���;��l}0~׭vY�NQ����]�j�wD�L�i������_.ל�'��BkK�J�xF��Q�ę��yO=�:��0U�Q�W�Ө��)!N���c�Z*ś�;
���De������N���?���۩��䝐L�w�9' p�Q�"Xz�w��U+?���������J��^,[�şe��ƀ������Y�[/���`�.�q�o��� ���j׾��N|�y��P2�CLQo�ͩ}��lA<i��[[���W��N:�7E�m������y�*[�}R�l�N��Z�a|�^#-��v�t{��{ )�o�"w��J}�D���b�"�0