XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~ ,L
�ߩw
�D�-99z&���I�l�q��yC4��wt�=]�/X����po��D��̴_��x�ҖQ�\�O��1��3�dd�^���!&����k%�K�.ʋ%���C��Y~��?��Aŗ��e �~�D'��ͣ4�7�C�Z�p����ZQ~%��ԉp�]^��WҌ��pClSyi�����#��5�)ٜ�[���>oR$M��S[T(�uR��y�J������΀T��<��\ڄ78ʇ w� ���J\������J���}��DdϞܶK��+�}^����~n�����|r�<���VS��*\�D�G� �f��y��?z �f�pJ��Yp���3�{�Z��|S�p{Z��^H=_�a���s��ހR�L����q�rB!�4���c#�B�M+u-�DZ�[7�.^�ρ{żB��`��`>(������W�K�7�>���Щa6H�_�@���x&�" +�O�y]W��D	�YSz�36r�O\�!�ָQ��?���e��X"�9�8&v#}�vk!��y2#ŚR`�eϋ���;Ejr֘�����dBt�݈��a�(�rPmCXfVz�ȷ�![�?M:�]��d	��b��PeP*�3�}usE��~+���_����r�<���E黋�3}�ɳKR�@�I��v5�峚XS��|�jY�s?r�0$&PK�Qc[rv�|�9�pҵ��w@"Jx>�H)O��p]͂i:��u|4��H�Uu���� 
��$4���=/XlxVHYEB    9d94    1590�:�!�"{ш�����r�H>?�P��+����ѨT�]�r ���B'�w'���f�y$��A�y����B�����ϓI� �i��Q4���-�.ad�\��C�e��.z3�;\�N�Q�F����mU�~|��@.���;Ui��+���2,���gM8�|I�jG���μ��'y�j�Ǵ�Y�����KXC�H������p$�����d�~�4����/�>~D�[M&G:�<v
<2c|���~��������'�Wg4����5t
��	�//
������Ҷ����NWIk-w_ۙ.t���$�6�6ޥ:��N��`']�iJX=�.^��&�7�J9��|h�^d���Cޯ��w����ί	�Q R����rב<L�7����y�k����Gl������{=Oc��LwF�����`�=��h�A�m����Z��M/�� ���X���j?�Ib�п�CC���J�<>8�.��Ot� )��i�6�W?���Swb�=��3�-n��k�R�B q����h�������ϸ"K�v�z8��Zj�	�N�$�բ^����*}��y�7t+21e�]]%ʙ��k4�l@��3R"2V�w��D?�N+K�g8Pb���sq&C7�d���ٱӟB��۹ N�Mq!�d1)����J�������/������\�M�G���tްVC˶o��zZ��3X�-VT�l
N��2]�N)r��L?�4�)(}3(p�]Ԇ�D�2Mb�����a�-�M7#!}�}��	�۠������4휬�>3�+g��E�e_�SL���n�'uv�}Э�bE0;j�k�1��p����̫���j��Vb�	��Zb]��<bch��?"�l���O�:h��5<n9�<��P��_���o�u0ZA��y���p���ZKe�OZW��@��{��Rd�Z�	~ԛU� ��X-����--t�*��!%�^C*Ke��S�0w��d�G0���_l�>"Cቶ��O7RD�:�iя��EJ~>t��R�
&�5��9V���*ִ0 �O�4���ə@�a�O�|�x���X�p�gП_.�`��F��q@��/ug I�񷰥��h Qӟ��+�K��}�4�2!ҐQs��,k7�|��UԞr|ha��s/��t��=�����ע<5����(w���2,�	����Ǌ�к�}Z���ͪ�/���2Y:Wl�/��A5���j�'N+2��8��a(��o�\6��&�� �KP���s�_2MJ�����SWz�d�o�u~dZ�[y�ɐ��.
�5΂���0�@��b��Zd]P��K��}>`8�F���G%SE��#����ld'h�gŊ�bj	[tgÐ\o�2����%�qm���(������@���f�ƕw-�7�CȘ��Fp�LFĠJpR5E�W1�l��9W�}yP���׆)�al�=�6���@Ix�o��r8A:��w�d��H�z=:�{^b��]#�V�u����)y��Ϗ�ll�w3#�0+H78c�J���܅J���Ab�[b[�%Q�\4�+Iz'9��T�JK�VY� �4�*�+4qu�s��҈6(k��RC���h�]K��I@.;�����F�W �[>���6��A��"����fE'��n{�ެ�`��� ZNĚ=�� 6�rc�}z�ٝ���pu!dh|���^�U��}��"�g�na�	����N����"����i��v��-
��^t�Lvnc���kb���MJ�p�����>[_ҟ�X"&��@<�^�N��0�s�Q��S�x�b
��ki�����K����YY�p�	���we��]z)Z�,@,�5dp���R�j �[ ^��6�z����,��Ƚ�JB$(~c����Q����Z)ӫ��X�r$hʌ���ǘ_�Z���;�����!C��$�/�QJE7}v�,��4���tq��33C�oEb��B�.���V)�}�镕�=V�CE5Ě�d��'L�/�E"'=Η}gsU�GV$�(���|��A~ �]��=>�0���)��~y¯$,�o{��'ЦLJN_�"#�	���\���xkҴg�W���ݎpO;��72�ٷ�?��/v��2�Քi�[3&� �C���)�-�𵘩�Ce�{��S%�q��,��H������R��֨�2�j��;)U�U�#Φ�s=������d���&@&�C��l���T����-�Շ�n
�5ٶTrAw���ړ�c��d�<�;f'�3�u���6����(z)���7J�W��;P�A���h�E���!C����<K8���W�xZ�4T 6m5�vn�M�+/���]`)U[� _�V��wCX�C�Q�>�a�Һn3�6�}y�tYc��>T��8��i�K��%���>
�VK� A�����D�O��pq���˅��'��1O�� �ob\4�8�nLf�0�sa�?���}VhLO�;'�c��2+�}H>�a7a�ڵ��C�p���Uw{�_,O��?��*ʤ�)�I�uF���̋���n�>���Q��ܗ?�;J�+�����}�4fQt���[�H�[N����sl��u=4�U��Ŵ+�VP�)�]م�Л�T�y�%*WZ���yk����\�]��Э�p�-�uf�5ԇ���	�(o%�1����W��FI�hw�S����OR�:c{ۚqP7S ����A.�R��
�"�c���p��]|!pd1F#YQ���q�� �A/���J�"��o�S�D��p��=����~��18���?-'*\�Qp��X`�ϼ[��	�����;üb��!L��n�/�_s)']b�k^Aa��6 	���*�S�%��_y��B�ɣ>�h�-H�b=+d� ����[xk=����A@)|�F�I�7��^Y��B��;o�`�Ğcf�tzK7ܔ��K*ǐܖ+O3��ƍg�[[2�!jʙ�zI醱tӶ�9}������?[��m��2���`Y�� ��1��l�y�]2�6���e�u����%���N�E�g��v���
p�kG����N)�V>���2� a�t!�
�����$�\��^���y�ɶ\_��U>��� l�61��l�X�љ�l!SL�*�qr�v�7?�b�Q%��O�����؆�G��D�o����
V�V	�h]���d����j��7 �*��`�|r����)��B�����^�w���>�Zc�e���9�A��5��F�ٻ�P��!k�Y�*3T�A��l�$"�H�QG��"a���e>ܨ�̙�^���f'����-��rJ�K�$��mIb.Gj#&A�-�P:����l�Q������h��l��I��������#��2���;h8P��l�`�����1(���F��"i�!]T�8�Z�i~尢Iz����X��q��s�$a����5������uhׇu��l��U$eb�X�&���J���J[����P%h�����A��Jg�m���;v����ݻygbW�����=<ãOo���~�����CS���4�A��ν�M�S.��&�=�N����6�j��St���Y�Hnl?�f��r�Ebw%����P�d:���ƹ�\#�YVq�[@
�f^�Y����e����;�9fG�ޫ���:����{\̯�۪ŗpI�ic[����N��ȁ��7,�Pvzp,r�oB=��mX�Rd��T�eⷱ���<;��>��Q.���s����+��J8��H$��@a ����w�MH�f���tkB��O��G�aQ5��1���tʅNV�S��{�e|�G�R銉�E�\�����v��~�xt�UH�q_,]6�D�`��q�a�\�r�1�%������~T��R�
�{ �6BP5�ja�{RWSz[�풽涰����:U��[Ɣ/�v�ǿw�W�H��-�q�1^7A�;�^��'e��5��C=_�u|t�;���� �h���6[�#�G��	-Aa$D��zKx�l�J+vv��>�([���r���*��XM�Ĭ�ڷ.≰�V��(_R� ���xm�k~����r��$9�1r�<����] _��=̗����K`-����3�A����"R�Y��Vm�N-����^�Dk��_븞mˎ��]���v]��ko�����d	���ph�<�+Z#ώ�g y��?Uf%�$낋�|r܅I)��)'�q����䖸8��ΨZ����u&�����Br]��ɫ^sQ��?Dut}��3ծ�Z���.�K�-!�*��V�/B�#�$������l�@�� E����L?{�N���N�\�5�wg��Db��y;.ο�"���M$��6�1��`~��
�CeO��Ѳ�]��.8�x���sTrQ�N$���� 6vؑ#����OdS���Ƶ�mU�D\����<�r�*��u~O� ���`×}筆Ԫ G�����a�#�PƓ�0�T��W�(^!���x����ׂ����ߢ=h�Q2�q�,�[��ջ��~�b�*�ۉ1�*�2t��Fh-�#�Z?Pp|Ћ�)�Kkמk@�TM�Kb��.8w�=���&^��Q���{
�s�乍���2� �H]ktA���_�cҮ4�K܀9���.aG=Ӱ.��s���ͯ�S0�rw�2�� ��T�	�u�L�&�sK��b=��N�~u��xJ^<��2#�9�U~�۫�\t��K��q�3��n�;���͵Cn�*Gb,""�Mm���\%�3$y�d��9<'��~�8�w�\��5��9Ó`9����ejY�ұe�F�ڗ�m��N�yr)�i�8̦p�	wզ-�u��G5����[?Uس'Kく��3![�E�����4s�t�����Q5�C�t���%F��2,����JHo��cd�D��k��dG�u]�:�꤆=�9��~D�$��m���~i�|m��dƓ  �7��V����\v��jU�g�͘�M�>̓��$�X�Uܫ�(�HM�/�* C$N9N&��8(�e�FlH�X%��I�*6F���ܷ�@c�@��AMIg�h Ɍ�<�}/���������KךCU�Z*��0�RjMv�1Ґ}Y�a��d�����e��SL�+>٢�c���"�E!^��l��������I��8>	/��b,���t�ͬ��HU�f���>$�xe�WL�,!�i�t���CT�E�|��No��\P|���6���<@�E5���9��K�Q�2"���u�h�EL�i��ai&%�$umݰ�<�	(y��L�P�K�U��
��ξƚ��@� b��"Q�y�,@��+4������!(X�$���:��
�g�2ؤC�B\�F/���Z���ư�����4��F�d��Cl��h�m��fa�V