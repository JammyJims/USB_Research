XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� 6#V�V+�9��>�r虚��7^�|��63>�Wt
��OX����'
T�(�6�G�L������r*��D/��e*�&-C�\1x�����j���("'L�@�rw���;���%d��y�!�{�bi���Q㊆����Pl0�6�Z�������k�K��
�[D����3g��:hp���݅;�-7�yJ�G��n�[K�R`_�0�fE�LۖR�gh�A���l{��[��
��w����;�d����vvB�T��W�_A��"!R���]ͺF�_�	�0H��@?��B��N�j"�D:��<?���6�r��!����x����d�^yVMP��T	�.���Q@��|�sN�+#[=���b�@Ɏc�Q�}�i��|K?Q6�cy�$�(�Nezg�)iT�� ��s��ǞZai��m���l��ÃV���	z�` �a}�^��%��b�a땙�q�K���zZ\����~��ڽ�f��gTj�\�C�Ϋ�%yz"<a�����#?���g����c%ݫ�u����O.T�u�M�_|�,:�V�s�4�ȸ[Z�V������铩r��5d��
�Q_�6��pY�!P�}��|�3W�>:E�����w�R��|�ئ,p����O�\c��O���pj�>��]�"C��+7�wR����;�U�Q �+���������AW�p�`L�:0�M_.��"@x�>H<�u�۳p�*[�I��'����W�߻��]h�qfl�&'�XlxVHYEB    9368    1370It/�n��̸�b�� �l4m�������dyˆ�E�������Pp/�������M'�H��N����:�'ܦ�#��е��Ԫ�f��/�x:�B�^^6�����("c:�? 8Z�H�T'~����̬���N�Q �j�ބ��1���ws���~����-���',�3P���}~6Y��/|�$V�N�� �2����pClw_G,B�Y�=��vG6�G;U��Z�-��!`}�N��jb´o��j��Oڝ4����LQ�~�綡�mCk�p��6yE6�݀���3�Ȗ�QE��%�������[��9���:o��%Xy�r��@oCo����TRr��Q������� W��˄�5x�H>�k���t���K��Y�Y�N�w=�������"�z�3`t_�)j��z���k(�7>u�-B����^�(w���̍��r�a�95��aEă��;xJF�'t����@j��}`#��u���IMМ����3��`���m��/� f�qfI��,�>I�NщX`ZKa2�jk�z\��/gsG��߾�����0�ξ����F����hP���]�)�<��t1ܪ>�2)|�uo�;͠1�twB;����DՑ�A^��>�}�����D���N��t�f��,����5�P��<���M	���>8P���X]�%{�r�h��_l��?2���I֩�4OMߊ���{f:�@vɾW�`V�&�>m]�2�J!���XBM!�����_7���?��t�~�ɮ��]r2�(>���&�>�	_b����iqO�opZ����q��\��C��8T׀��z�ŧP��I �[�b�Q��	�����q�W0zq��!{�SO)2�J}Wĩ=�qܠ�J��AǝD�V@���7�f���l��q�)	��-i%�hf� �ȏَ����5�'�A�F��*��z�󇙥@M�^�4�#^0R�X7za~(:�q����%�I�.�7���}2P!�Q�t7�$/��?�M���{d}���/��`o���^�%[�81a�fM�S�NE�e${MA����4ӡ�h#PjP� �aܳv/�T3�������[Դ���>f�푗/��R�u��Ư�c)�=}[d����o�yXj�7�JCR�=��F��_5�nѷ�x�5��ë5[{EN�w�؜�cN�t�"��h]��=�S�Å;�| R��O=�<�G��7" �-m�Y��ءL�hV�I�B�h��jz�����aŖ�&��2��n��Z������[���)>j#�FQ+�S����o�q�N�.����:gb|�!���tZ����ј{P�'h_M���f'K5�H5��7D��Ш$�O�Q�A�"���2��B�myHyo�	�s�����z�62XB
�@'9���q�t�a�)���kG����i�h$�y
���l��Z��%V�x91h\ц7
���M�o�,@�YqfeVH�h	��K*a�!vO�*��)�_U@��Ǫg��f��Siq����Q�EK�m�b�3�t�V ������!����I[���^�o�A7�EqE<[ng�����$��NO���Zh,�V��
 ���;qC��S�)���ew���Zr�����F3e���x�Q�4�*��v��D�P]�.J�<2�� ,܅�o�Գ!Ԅ�\Įv�R��5�b7�T��C���{��)��7/�w��sj���E���ZaȊ�����v�)_�{Į%Z�=���uR���]�1	~��"|�^6ޜ�1HФeKV1\�Y� �$�� V��p�����6���Z�IҸ���k)K�tms���T���/XnHT��W=��r��a��g�<�d,�u\
����W5�Q.Ͱ@:]����y޾b���D��73�ĚZ�����ɶ������QK�����(W�ꠊ�����@�ȬOmӐ�V4t���\d�@��#fidH����|n�r70��*gس.�N��?�/G3Xz����T��K�����c`k�bsA�O�����ȸ���8 �wU�KockR��6�S�� ����S{w��i��ɀO%��rTy�Z���e�z�P��� 1v�>DC ��I��W��:�
��1[��2��C��C�G*�x^�u_��'	��%9ֳf25T<��������6-0��b(��c�R)��YϚ���?ٌ��5�����;9��룏z�N9�a���v�SoP�-@�2�E>��rYs�x5��M�̷dz��/���ф7����	bV �t����1��E(���^�ּ��a�x�k U)���"Hm��
p�":�by>��5�
ft8�:8�'�K���y�k
�Os�$_�ቜ3�vB��(��[�{i���u�z�9�nѢe��џ;4�[i�[F(�����F#�\�5Q��Bgk���KP�[B�N�yIL�s�I��j���Y�k$°M�9�(��>����E��Ϧ3���gNCo�E7���;�(�*"Κ��
�	�Ŷx���pXM,�R�ӳ'��5� ]����e���U�FT�G�||�N�yCu���bTc�r©��E�U�r;��@�H�!�Za���n]�Y�+EA��"��Ex�v���/,!�����X	s�'�����y{u�\T�-��uݡdI�)O1�V���a1�(w�h��O�4��T����GsK-ei�'�Bb߀q�@7	���u��8�QZ�?,�^b��i�.o�;�WC̚��Q�?�
��*��n��p5tJ#m@Vh�И3�M�X��9�&~4(|:��;	L��T�:U~>� 7@�[飷�:�q�6�aY �*�Է�+�?�0��E��'>��i����!wG.�]%`��T�u4Ri[�M6�/+����Cʾ�!��� ]���u���܍)x:��"q��YxR�,�i���P�f0O�z=��u��"�����ئV_?�\��!3)�������5G1�G����t�+
����������3}���qwXkW�rϧ�]��)�25ڮ����9Ŝ�H�G��UZ�Z���ܚi���X�8ޠ�#A���O?�DXA��,��Ov�OX(M���a�~�g;	�ܢs"�:)
�P�A�O��0A�=$� д\j�2C�0y(�l����WaO�:���k�������
+�h���PJ~
��{�{����<~@��6�G~J�����9st���Ў=U���}(�5g׋&?�"��=̑��/�P���^���>��v��n�h�n>�{���S`���7�>L��A�Ko�Y�QC���j5/÷V��E���џY��4�ћ�:�*Q ���F�?/Wp��{�Iz��I�2.��{�g������������H˂�q���b����
@��״QK�Ŵ��4?��:�n��,�+S�*�f����!�� ~?T���A� �m���[�~���������fe]Nݣ��$���e"�_��wlnӔ@��b��yf��ٖ����4�����1�	��ڋq�kO�E3�����>m�2p��D>�m���9gB�W�=d�f����J����	�4������L����b��G�Yqi��R�>ޚ ɥ��a__�Xu��&�_7+����n��]w������ [�ν<��B2�G���u+	 �?�隁���W����0x�h�v��(�%�?��@��\Q� :���Fq��-�s�^�,���,d�k�n�7��#.�-{����}��]��UUFL�OgC�_���5�N���4?�i��`b	���u�8
 ��"�1�p)I>懻�$N��Ћ䕍�� �~�/�UaBY��/��"B�1Ƌ��w��~��Xh�ù�%c��������d�1����3�R�LG������/X�"��b�<�rJ��ݹD�Am�N�5C�@�L� y�o�3��p
�� MKѸ�'BK_/b�!2i=���d��]�����0�M��iL���Ҝ�lWJ1|3�vP�}n~��G;�|� :>"�H�}�쐕�^���j~>
ʼ@Ԏ��0�|@�36f�?�m�T���8s�K���{_�yi�gM{j�n�y����5C�,����L�m��� �$�[�e�|��/��V��d6��#S?�3�6��刯A	Uk=�NbK��/B�#B2�uQ����U'�?Su�ҥ��_��5�N�J�jm	3�ju������x2˧��P�8�(Np�.W��?�7�:Fc���
Dm�B�������DP����� �q��,�������y�����O�c�*%<��\�R]�N�����y 3Tr~���L���2�8G� ol��N+�i�G��|W��+{[�>�r$g^ F>��z�U�������]������b�c�I��&r?��#����_J1W[$/���7k�9�\mB H�����1�YYm�	z�G�K��^�/u���mC1��9�y��]��,�(�9�}�?Y֣8���N'|�F����0+�d�4Vw&A�ǥhN�mFF1=�$��	�'K�(�O�3F��ê�1�SX��6_v��3��ra1Ÿ�.��r���u]�ke�%��x�?b�D�U� ���?<jT_E���Z��U#2	���[���k�*T({@�a���п�C�������ѯ�&�@��
����=y�L4q�t��)&H���8�Te��o��e.hw����C�Ƒ���lm�?!0|�5�Y�H���.��6EfH�-����Q�Q�*��A.��6�"H���q��<����w��Y�CD$x ,~��T�|C���3����B��9"�p�;�Q;`ˇ���贁�0���wܠ�.ț��@)�� ����/�sH����UZ0;�85�؇s�%y��� �n�4�=�5��%��ȟ�