XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c+0�e_3=��a+/ �Pl%0.�?8/��m�T��~Jǉu|#ơ2�3�]��e��;,� 4Ӕ�0�%T�(���UX�&={�%��|�aK�c}�tǗ$LP�x�e���tVs_=��aZ����ǝkB�^��Q�
�t!>����
@Wr�2px1L����LQ��ʏl:�-a��	��w�k��� w�;��v,����mS�x����������
��UЦ�Ը�l��h���H$2����S�P�������2��g0���?�PX�]	4�N[��^	E$��~ Hv�cT\��{n�P4"h���<2b���EP��I�Bԫ��B:�ۇ�6ŤȮ;,�)yEb��7�ƞ�� �>�o��O�tc���LDH����六/�����M�_-��S��`+Z"��=�VK��L�1�x�#����&�ݖ۾�|�S���U���"	�β�*�-���bJ�ĥ;��7��X�T���\`0��-�j�`]���??lj�l=�aUw��R�˘*��N��ut6�5�	)DH�6_g1�xzY������[�V�̩>
4<�>�A7Qz���T�p���R_���ӄ���tq�R��5RR�߭����T΋n!EV	;���fa�U���FΤ����jK��~ ;/q� �x�����'�Nx�"��z�k_�iо�V,��v��ߥ
�H�H~,�����!�@3R{���J�{Ϥr5�-������OP:�/�ΕyA�����jNA��TXlxVHYEB     bd2     5e0��v�	�� ��3:��U�O��L
E�j��߹2����A�@+lۀf��Sv��L^�yc|��`&��x9n�� �AH�C5=Q��R�T���qRE=LO�>��ҝ�k?wk���o���h�m�0 Eכ���4E�;�!�	�R����r_:����dw� �1�_j�T��e.�s�B�^�G�^(���:�\�l�*��C��2���ڜ���t1������؀�R�iXN���O.�j�t�ּ��֧���k��eI1��kj�^�0�bp�c����,Ȑ�;�T���0�)���N���
�S9���0�`j�2�mX�80�ξn��Z颐�\���u�ZVFd��!��9�� ���|ԏ�d��Bץ
�Ci�f߉�� $s��yɥ�N�;��{��t�Nx��Y���XBI������W��߃�����-ow�����H#|ٔ�.�7�����/n�ck���l���d��V��Ӧ�! �����%^�o��P�G�rbr�4Q[N�_.�7�����Fl(q���ɍ��f��n#:����� ��l�o-��|�5K�ک�X
�t߱�I���o��j�s��|Y���l��󤩌�!�7�1�_=�EA5FrQ�\�a��#��3��U�C�p~g�P���ǟ�2�!�n�s�C�^&�|e�oXϚ���/�K�z�'�E�J��"����f�	�cBa�x����b��'��Nɒ)����שЅ�A�=��d�zHȼ���J((��}���xxKT�4���	�mv���]�<�z&#m�M&L�2��h�!쫔6g�L:�i�s,�G�a���V�w�����K���9"p�*�6:�j��}U$�]�r"�� )��~_�Ikl~��y�.?/*�����Z[�)CyP�0�T�De�'��&��Z�7�[Q�{�ٿq�.��������뚰'+8�/������6�,N�Ⱥ�3��8��c��H���nӜ�JGJD�����Su���,'%�ؗA ���T�*�>���y{�������r�w�ON\G�u�=�
z8��!�vT�n]fS���K�vD�n.�H6?����)+�Q����0sEU�hX T�^�&���T�[^�c��-f(;�%Z������ye��w�S���4M"h����%8��A'�0��~�忢3y�E)���B>5	Ci6��$�������$F	��&����A����m��.�L7�8^�7t*�;���K��ty혫(x��%'�F��J._]E_e���K�"�M�9qrӓ싪]�a\��M.1�rF�j�+3�Qrj����w��`�T�H�4c$ba�K���4�;�:]^!��j�g�׃)���l��Ǡ�-��(Ѯ �p�®GCm��&j�zk�YɥA�U��ιDPO1�c�'�����,X�/:YUɾ쓫<�30���u����/p�·���oc��KbV_��)����kW0T���X�A>Q{�c�W�