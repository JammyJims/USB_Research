XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O
FHg��o m����왚`[���FG���p�	Um3�2�FO�F[��$;��Avu��n���ѰT�eJš�$��3�uH^�l�� @g�|���L�.y%S�_��^:[�]�c��_����w�>{�W.�S��&�6�\�f�鸴ų7�S��u�®��J�[����ޞ�p{��-?&����B7!��W.Q-y�d�$mXD�#|	�F���;1��xzOW=�ƍB]1>�����-�����nO�z���W2�@��<�:�����%��j�+��#��V4��H�Jj�z<+d1�𫦛i�)��+�H�x��~f/M�7{N�2|��;��;�0�d��E5�X�� ��A�5(-w7/�ᑹ��7�:ڛ{��}$4��={~���؅|��͝��QM����'4�L(0��s�9հ��I�}]�e����r�0m��w[�~��Y)`p�X�qQD�UF�g�����XM���">��X�ݞ��-�*��p�.���`F�׿Lzg�4~�MAK��� ֪�'F����B"��� `j�/c�;P@�smL�.[X��6�*o�Y��w�tJ%�o���߷	w��4�������Mv�͡��%��%���E�gm�'���.1�05b�^��2����\���]Uu;�x�� O����ѫ_��LK����|�v�܋u�h�!1�ŨQ �}�]���\�|�� h���)�-F�y�e���qn��!��w�:���-�+hR���U����6�˸N�=��KQXlxVHYEB    fa00    2360_]�]ۆ��{�zOǢ�cd�)`���ϟ�s�3�q���P�̩��F���l��5���Ŕ�� ���W����p�h 3�ŭ#)/��]�L�e89�^�g�R����<^+)�;9|^�����',R���]�H�T�ȵfx�E�|��:*�f�1b�� Ӿ�Mk��yG>��Tu��!��ϧ~,J|q,�m��n���g��X��Ē�,;��TeB�V�$�i���_�5��ӋT��N�ܞ31��$�D7z��w�m��@ls��(7`@�w0�ʃN�G��]����^j�H���%��J>�ę�ɋ�x�3��k�;C���y��������Dr�=��1�IYk��1����E)��O}I�]+M7{�	%Ú[p].�
6F�9? ~ ���
hضm1��sm�N]�Gb�L�3J$귧~��^H+?;�/��vȝ�d��a�qj�)��5ߛ�������[8OY�B�z+MlG���!w>��JAO^G�_[��I;5C�A���[�#�}��N�o3&��/������R��
�<,�3I��OB<M���g��H��v�����{
ժXth����+���M�3K�$l6�׈h���wF�3_�~�޲�ê�ÿ��B��C���l��O��=��J��y �\�$�S�ͻx��k'���*=�d�G�D Տ���hc�=MwP�rz�]��KZ��]>ǆ2[˩o��;c����B�ceMuW��*q�r�V|��h�`�oy8����$�{)�!��b�� �g7��P��-��5�vN��&e5b���QF���ux� \V?�O3�E�ŋ�����^�cG_āT4v���mL^���@x�֥�a��HxA+)��E��$[��@a����Q%t�)xO�m�p,�"�T��謌q�o7��N	��]pUn� Y����L�T�A�*�	�J�O�ʷe��a�C^I��l9Yh9;�Ҳ pc�l�K#���>W��c�	$�x�)FF���S�j�&?�v�g(���_×Z���*��S.udlo�Z�R�������_�������:���a8�Xcw.�h}��X�z�ɍ�	����$G90��Y���b
���Q��RI��۟�,�,6!�l	�|��b�c'%��.�З�{�2:���o�C\��yIj�ϐ��髮'
+�?���+�����p��N60���i�o�W��s����#�/�1���:�SFLS!JJ缩~���S�v�f��s��B.�����SK^��v���<T�ɺ+W�	�ƣ�vy��U��cX�?��l�ey	11o����A hftd<&b��5R59��l}�ǖgT��d4M���WA�_	�>"a�+D-߭�e_�x=c` �D1�����P�<7t�J����s�"J��M�B��Mr��[R@�h�M��1*���My����J�����U�
~Y��|�C�¤�K_���cOx_p��[�B�%�|��=rKD��s��#��u�ں+SdGV�d
�֯c���io-c���>d�0�:��(P��b������J�d������c[sb��W)�U��@<ĪW?��Z��t�mL|��E�F�5U<m>��7����)
u͟���6/ ���b���� �K��B��"��-��N�F����pec��v��E��M�Wm�w��Gm�ܙ�=o�ֱ1'�<A����zu
��ʷs
I΀ۉ� 	�Q���T3�r&�N��||HO�v"���Q��� �zIa���Dd���� �iA�{�L��m��*W��r ��9����lN�K��!tv�̔O�%���y9?!�}r�ŐFK/��ǆ�{(���]m�\���n%I����lQEb�y����}nP�9�[�-1b}�v���U<4R�F'�^�:�%+
[I-�:���]/�g=঻'B&=x�o��3�U:X}��G���ޤC0��X`*�MK���Y1S�6�t�Η����+�c2��m�`Ǽa5����W(��vY'3"�=T�(�+֡Q���W
��}�z_+ö�����s�4�� �B@����^�aRB)Ew����)�$6���!Ex �_�的�̑��_����%�jDm��u*3�-\�~:`D�k�CI���ꈔ�ط#��oUj��jG���/
W��S����8|i���kp�3άD~5��C�󒃓��P���F3���n���0��x={_���SW<�͏��	VJ\�֏M#�P�s��X��/:5��T�l��*�Nܱ�H�X'�f	E�3�F{�W�Ya\���W�k?�D-�Χ���Van��%r�\)���'�Ƃa����+�I@ڨ��r�FF�g�h���OPd�����v��q[Ĥf��L�aWW������<@̩#��W 
�uh:ٟ��aѭ��6���@h��
!�A�w)\w�������c�
˒҄�'G��޴gH -�Y�w���6�^��w�	��C��1GcKo�y�If����b��7p����DJ㞹��i�Ģ&���U�pk��Aj������fƂ��sO	�܊.�x�ުzvC��ӓ�$��f#-���pN����d�����	��e��OZ��?��4K�]�Г-mK�u5����ZR����Å?��]�S�Җ�K����i{~���3��(�g���q8}�u�H >O[}���g궉\��8��p�\��Ԟ�FY�x�]U*Z(��V%9NC����H���c�#�G�J�Y'?����[#����f�{������Ά=��G.�<�������oh��Z*���ߨT�U��ݎ�C���6Wj:]W�E<�H�˰4�Gh��}��B�R�}��ɛT%�4*RDz�G��}s���1w��wS�E͌�z%0y�����#���I9�����9X�]^�7�`����@�#1��#2T�Y^?�����ī,����W���YHb�:D�a:	�0囦:���E:�զ�{��P{z�O��WH�������n%~p�O;�E�#� 18f[[�� @!�
�Y��&���rk5]���ku)z��6��?�>�5r�á��5c�Ǳo�8���Jb�H��ϱ�*E]`D��ڂ��_���G�r��A�&�,��ɏ�X1~����w������/4�������P�����a4� ����X�nw5�B.vRp���;Pk��B�%+��4+'����oh��������1[d�h"ۧI?~+���0���aL~�&���u�uD����|臘� ���1g��3D�VU�����R�d����)00���(fL�W�cF�Q����۝�0�_ K.�#A��,��Sk�3�"�?M
fB�|��2�x׬��e�l?�����?s֧�߯���SqZӌ0�$��V53�z���6�@
�ڒ٣�����hXN1��R�"� U��|h�I9-4�g�Ki��o5��(��g�?�ĹM=�BgjD�9�P%�Xx�w.j��v�ܯ��ߪ�����CK����_\9o .�92Jj�����Dl]-������=Yw�'�\.��\�{w���z�IW��ĈVejY=y�Q~c3f�e��b~�����}̔ZZ�TM��%~z|j��u�aj�x��iFC���䎵�YO���hK�W���P�Of�VI��^ɵ�3�n����|��K/��tL!�w-ѥ&Ð.��B͠c���ӭ�ė�6�x_g��mD�U�h�/j��"m�ޏTv���~�a��|0]���T0�e��?D���]��8��+��aiXk��[�O���Z��T(�c��=�D��\XH�
X�Jf�{�ا�����/����f� ���+�M�E��7	_�@$��ě���o�(�F�%[Yy�����u�JN����{;4��ڄ�p�83Y�_��W�^�N����sÉz��=�/���d��_�m��)��E\���im	��/��1%ߥ�� �K�M*��u޵�*?�G=�Z0E9�yn%em񰱜�+&��O�4�u�����3�)�z�j'�s޾�F��T��K���@��}���7A>���&�XH������7�p;1|Ħ;&���Ԏ�[�)_��n��!���GR?�0��:����9N���KJ=@���������\�ΧKm�|��(B���{��Ǿ8g�1k��(=7���M�3�G�:;�
�eһ��E��p�^w*���}ھ���1��I������P:^y6W����*�FB�0{j�P��{l�Q�߮�"̺���h<�0�;�x�氱����T�BJ"������t{��r�J����n��x/a�w�h�ԣT�Hi�AŞL@���f�$Ӏ#D��CN�	Y��9��~@_}�F�Q���B��9>���3��v����V&�j�I��L�Ko�t�� �n��x�shÞM�%�x�h$qsw�~S��2$5�ћ���5��U�`�����6M��J��]ю�N �hf}I� ����.V�{�Id�Q��z��/������zĮ}'Ǯ�7�0���E��v�����+QDu���|�zN�jX�E/�~\� F΁���"�����<��GJzk���,ƍK�M����x��lTF�O���T�6�AE�����Խ�ԍ�Ȼ���@�,&fT�����ǯں��v�O)N��6�o���߬|%v3��k�w�+�nzށ9��I:i5��?��5<���t,ǐN�������Gș��$l�� �ɬt����N���ls�x�O󂴖���U�&wD�H8�)7��������ƺ~��nf����@(��]ա�QY=C�H-q-,T��i�	)wB1�@��d_&�_X��/O	�&���) pV��	&�0O~?�P`s��PmVN����^������,���%�i�14V�Ȍ�����)�"�ߞ�{�]� ^	�
���.�����,��7�K8�/�\τ����`B�2{��CnM�f�uم�YD?LNf&ƃ�wSpA75Q|6���C�.���{m�r����s�'�LE����9߳�ԱBCx&�����f�iIq�9����}Ǩ̻L�zӱ�N�n=g�
/��tQ�}Q_��jv�b�M�����i�����X�h5|9��e�j�R
Tҥ�w�t�O��Ƃ �~�X���>�1&p�|��E-ޅ��8H/�x�T��\{��͸���[����~@��n����]�y�Y�5��m�k��ưp��U�6h�h���C�.��q�i��.1"1&�^�@Y#�!5u�@6�P������`?��k��e/~c:\w!w��h�[&)��P�B�����jL��Z%ڢ�ߢ�ř��>��;?�#�0Ý��X��������B�^������i�R
f���&��'S���*0}�r�^D�s���"�	����$I6j������e"��E�$�S�sIw�����'(��Y
o�ȧ�� i�����\���QO�E�]�����=g�x��~���iHĽ�h)C��:��Q��L}�[B��]rh���}+㴤���T��Qgń����� x��-ou;�u~�ZܒC�o�͚����(��z�0�,�� \���u��Y�ߙ����S��S)���W_ϐ�v�F�	��gT�̣OV���O߳,uk��y#蕬m_�U��$Vw���>ķ�=��6��2�&�
�A��:T�Tj���I/E��}�E����;�U�v�_�>��N"��{M�'"!
�F�� >��_u�Ț	v�yuo�u0?�7�Ҩ�;[B�'���_�o<e�;2�� l���ΫK��,ϥ���6���桁��x�+�-����񶰘��zT .2��z��9���Oi� ��5�2nʢ܂/�r"s8����z;ζ�1�:�j	c��C����Ơ����f�1�L^l�K�6��Ͻ�����H�#s�ح����k��	�2��W&�=�>�o��m��*_�x�3b�	�@�����l��_���%ij;�6A+�ȟ>�PMZ�Y����%�O��Mz�*���G�89�ĥ�A
��Y�;�]�%[����|]��Cz>��]~V�a�%Ta�s���@�Y�R8m^Zn����+�o��M�DD*�"�l��-��s���FR}�Z��l�4���|'T�+ ���=qe:z�uu���.��.��]O��<���ӳv$)'��SYVS�u@���ʳg�@S~5�8�C�?="$��R�����ڈ+���w�3��1Ա�֐\�Rɴ�"��AHZB���B0P�[3T��co
��Rw����=2��L�=�H˻�wA�Qo_��GAo�oA��q��8��h/�g9I{�{�I�:�_�����o_o��ܓM�.l�{�o�=�Xm�<�3	 �L������M��B~���z����d���~��"R_(hlP-B��'R���L�@��O�`��<y6��ULNK��^Q\�ɭʅ6�K�fv�O��o�{��h9rY-Nb?"|;��9@�8P�����9	Pذ�k'aZ�E�����ٓ��V���{PN�A #VS%��q��)��EU���&1�dwZr �����pe1GU3�i��}"
6鈁�i�&�urԕ��\ E�I%tFV��2�T*���2�P�mRc��O�q�F5D�ጶZ˾*����<�t��OT�e�g8pȾ���=rs�6j�����Wn���\�ʤ��@��<]��X��
���Q1v�I��R{���锲T��ʁ� ���DlgJ��+Z����i��hw�Z����(1sR��:Tt�^Yt��`{=�E ���S�������d��A���H8G����4+�S�v\X���//�HLݜdɟ%�oф�!X|�3(�<������+��YI���O�����s�k�Kb*'�՞�HMEӴ�١�"���*�`�Z��#�2�td}L�z|��o��a!(8�65��g9q3����՗0�8���+&4�e[E"��3@�vRX�`e�f. ��!�L�֍�2xs^鵆6���8��L�5"�E�.T�5���-9\zQ/|Z6ے�*���q0��!E�0;K5�}����6����l��q�4�s��
��mIa�("0��]�n�bvzNkV���F��p���u}�	ү�5��T�ȁ��&�c	��bPСA)�a�ztS�	���bT5DK==i�-�ϝ+��a�E���_y'��_E��)�l?�Xk�Kh�M�z���r�]��I6.qu	��Z��{�Fg)�����%�
��lv��9��M���k�;�`֬�h��O{�
<0P0��%���������g��� ����v�4i��T
�v�v_Ѩ�/��7
������~Y��ڜ���6�n/<�E�z#��%MR�KG���	û�]\�`�%6aB��N{�R&Kx����͓cÊ��>Y�M������ l���8�0p-�1ΘpN�5�c��+Ra	}�N��@�4_�^�;/��V��j�F�rf	)������ݤQ: B�z5ʃ�	<[S��G���P�g{�d�w_~"a��h�5�v�F�� i'�� ��Xb���5��R�J�m���Mo��Z_�sd�x����=����L��n��UBs:W%D_*ӈ�������O���A0K=�a4�4��w������R/�]CU�����������Orp�kѫ&����1y.�8��ìkT��@��;�A9>������?/o�"D1��[�w���:l���:������dڀZ����!�aXC��=!�M�/S���48�����3�Aہ�v""��ҀȢ�!:�6���0���3:�ޙ������wZڤ����g	�w�Ы�� �bG������;L`x3��N�ײu�qn��HڂAv��r_P���ꌣ�8zT6�PQ�O#�j�0'*���~�x�s�xP���;�hզ޿<��Z�*�8a�B��F�!aLk'����t�5V�Ώ����6Xv���x{�����2�*�{���	����G!�Ё��x�/5���.�����O3E���-#
Yԍ�U��]7��0;�Ѧc�p>c&Q��e�����l� �G�1Y�:"�zo��n%"�(�ň�5C��z�9. 2�q���-�o�
���h�]2�"�O=��l�GU֐È�G�fe����|ڑ�S���	A�T�X�N�wX�ڗ��#
�z�I�B�.�/-�;��@�!Y1�+�:��C�z��'b$L�z��3��-.�Ƒ�6nC���,n9{�%T�^KtT�>�o(�*����BeQ�8Qc���4��.K��#��1�u�1��75�B� �m�8<;9��k$A��K;V����5?r��K��6U�92y��	�\�in��#������j�W���##�ִ����ƘߪWTM/"1����(�`�ܜ��� `���K%����OʮF�ߔ�����%���������v�N�'�������:�]z��ѧ�dU�7�t�~g'c���Pc8	)U���}�
�pkQڢ�0�],�����ó�|�/TK�J����ިD��=c�7�w�g�T��L��Oe&�ҩ��?kW��?O�~����CPNk��ň�^Y4	S[�����"ֵ"�а�'/SK]�d>���;�i���;Cs(��~����I�ը�?���<eBҁ8�e�!���f.��@BOD,$�4�o3Q/p�Z���|qK�aosZ��8US�'3���R/�W�q��������51fQY#y	H0�����^�÷��$�8�m��Cו>B��6.bΜ<����q`+�9��b��_	@�9���H<X��Ӹ���՘�3 ��3YQ~��J
)�p����,;�~���롂����{�ᐽs2���z�lv����z���:�=���\.�ႆ�>
o�XlxVHYEB     960     220+LGЈݫ��Q�@X$w��>ɝ��"����vB3k�J��D��	-��H+���/��چ[W�l�p5g)�g���xGl
���l��o���K|�O`*::�u%��L�4��n��{�H'("h���sHE|�rR�ov��#��]ǲm�C�z���Ų��	��Ϗ2���0��LȤP�j�A�YC�-#lTN�BOz��"�W�|�oJo�G|����x�.�n��Xm�$�c��9Y!ϓ����@����R"t-����P�.��2�������4ݝ����[�e^��:�&OfB>I�̄��d�~ڂw7�j}�ꭴ�I�%�q.��i|�>C)����_Z|k�<X~ *]
i}m�@㈏#�o��]�����}L\5q�'���h��XfSz���}���Ur�`��PX���ak��`uә�1�-C&���Q6\N�l���>7	w���z�f;�r�U<�ѝ	�;���*{Q�5�(��fp)��Љ������Gߏ�������N�
T��