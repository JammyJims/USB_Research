XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����*����{���B�W��'�<˙`�L�~�DU��~��z��ж���3lb�Y�s+��;%�9z(�Vn�jhk§/������&�C���h� (�ࢂR�BLCE���Gߪ�J��Fy�^ʹ{�2�EXh����$Rv�F��b�|��Q7{U�c�C�C��X+gk�βܫ�����h��a���$��sT��L$4Cy��<bRUq����^��i�bi�cx�t�g|�fN��QD��`#���2�D�6#�FfԀܺ]�|<ΜH�=]�%�9R����eu-$`?b�'�N��`}����Y��(/l�<�wv�d�o�Ԭ�#1.��(9��Q�|���&�D<�Pu��m�%s�lgGS-���ø+�7��-��XU7�g��[���{Ȍ��IF=-��]{s�Gܨ�ʨٜ��;�S�d�d}f���;U��4�l�� ��-��h2}��>0����W{4������W�� z�3� ��v����mD�BA���[#Ğ�v�]f��qG%�%G��+������	�Vj�u�}}�餞���>�uk�D-��?�K�d�tl�#���c���-A�I�mڏ���Ą�h^�=��p�XWE�� \���|��9��/_o�3ζ�o�h����i���By��!W�&�Ǻ"�w2$�/�,�=+WXd'l�b��޸՚jY��7���^Yҫ5]�8�kY�e��ؗD2�ؠh�N���?t��˨�	��B�[�0����!���L5 �R���XlxVHYEB    b7af    2960�V''g礢s�k�^�p�!ۙ�a��}��A�'�T	�h�z�
��|��YV��ղ!��5�1�W�����>3�yW?$	L�0����Y(�,׳d��1S���"v�\1��������;���X���v�c�]�^�.��v�<���z�7�		��s��T�"�sE�������k��;�@[@		�Xb5�6��a�R>���i�|�<�'���E|����U��Z-a��EX�O1ȉ��Y������ݒopכN �@U����'��D����p�f���0��u& ���i�i�(��|����`?k���%��\ }��T�(:�����?�LO9�.�1�������&���� C'�&�T��h5�M	<~fS�v7�ѥ*uM���`�o�EJq{�v��50בm�ԉ�����ɤ:Y�c�,;O��6�����W� �1�kD�l�+0�&&i���`���{P�7����7DT*�I���k��Pc�d�D7�j�i�#�*u����c��ΐ?O�0p��J8��#��,���Q�7�=4��D���T7H�պ��;o>vi���-NhT˗�w�\|�\ Z�<�<���#��OUSq� ��L�ON�v�MF��"�y0T�4�A�e�(�z9�Z�º����T�H�"@������o	�K�?��AJ����\���]X	�ؖ�� 9�ez&'��ʹ@A���C-zYȮ5�B�CΎU�٤�j��K���(ڟ�K�����"%>�[�|V`x?v��y|�k*[���||�!�AoR�`�/og틎H�S���z�t"ͬ�}|�	e!q��p�)�tuH�p�b�W��C��B���85l q5��)pd@DЄq��o ��;jP"��X`$��F���,0��L��5��-��]�h��~�M�o^p�dC͎�ﾞ���D>+�0�'ǽ�!��}�o����͖�c|;�Z�pܧ>�5\�ܠ�/��]_��D"J&E+��Q�3�S�ֶ�¦o��ƾ���5��:*��������g�܂��᷶�{�O�4U����-�)����}j��G|�}��CȞ{hp��4�T[�9��������✶�Z�nA�%����-������F��>O�#�;b>����Y]yW� seh����˖Ve���̵�y����.lA\x8�Ďa{�Z�\��s�u����Nbк\}�/NI��i>Xg<�!��wJ(�v�t;!�Л���׺v����ѭ�s�/�R$�QG���X�B�u���a����=3}J����6]�!ED�~����,@��?����#v|UT0,wqPse�5I���4�J釶�>�I��!�W14���!B�'|(�(��%=n?���te�UoZ���NdZMW+Nq��~�⼫.�c�lK��jO1���I�[~�/�X��R[��o��)3�2B�gvN��x� �t�B�JA����c�y�Ed!0��:���[/:y����~�<�."	h�Bpe�rl�� C�bM����"����<x���98��#^�~�lܲ0 �ZD�xG���G�arډ�%��b"��0X���zW,���ĳZ�D�tXOD}��Fȥ2Yh9�
]�!���z"^��z{s����EQO}��>^?��Z;2��ܼ`,����)�a��E�Q#�n���k��l�fj�K�oj}o�_�[D���
��`��"��B���!�e6�V����6�;(ڍ�����*�o3|Ž������߯қλ�7Zp�S�S��f���M�.e�v%�ź��ҧey��ºa(,��NeD��K$����'̠Mj�]��6�iPwxm�# \��µƖ�N�e܏�5@�Aϓ��~T&D��C������8��iN��T�)،rZn�C��8�Rէ#.f?�ٞ��%>��/�CA�?�on���7HR�ٳ�R���d��x`+�L�Ydz�}�0�0���Z`�� �$�2��0je�-Qn��Z\0� ���U�(D�" Ef�|р������ܘ�)m�YP�99s����;��=G�I��<E*mhZO���q2�T^Ґ��)��{; ��Ir!��h�f�Sggo�K!Sp��*�+�Z��iҠ��uy�]=4BS�\��홋�ZD��8��	?�.�筫�-j��~V�S��Isa�\�j�G���B�� �%��j:A��K��c�Y�Ey)�sڙ��6D�ż�5� ˓<	��O�,3��f�`5,i,еP-c�[�V�攤�l"�N=�οw�c��n8儬�� ���j�K�a���	le")�����"�����lT��?���T��nc�&�<Z��6�k%ۗ�g�;ñr\���6���_A��.�i�Z3��Ʋ��5'aϺu��t��7b����IG�Ѝ�����3�,i�Ϯ�ӫ�=�YZ66�f�L��:M����z�4�Xҟ��tn/Ks3��bٺ�of��6/V���τ�n��{J�o��'P�S �����$9'`�x�W{͂��ɟ�9P����8 nP��E���iS_���ul��G;ef)���D����ݻ�x�l�Ɉ��4��~�C�!2�Hs�5�$!켃�܃���r�GBE�����$�u�"�$W&�|O��Y0|�����2_�Jo��,((�m2�s�P�%K���dh���1��|d�)qe1ǒ-�"��z�ȡ�Q#}:�X����ގ�C��k�Y]*E���a���J��WG����ڔ4L�.���W�-/0]z��>=}�Y�)w�����\��V�@�	wQ�Dk4;�a����lv��.>]��`c��ͫ�]�׌l��޶$�2g!���/�G�͂�w�������ڌ�'��ć���s������C��͵�X�z��+d�Y4�:�0�v�����̒97�6���w�&Zb����(|r�:��.�Ⱥ��~,c�_�Qڙ/�t�,���������(~ջ(GV��#͌ˇ{���q���;���_j�.xJe�g����}�!��qu�q%�U�m>���D�AG�!1��S����d5~�F��H�9Gm� ���'��K3x�&�s�#Z�Ԗ����,����WZ��%��	���"2��2av����g*��Q�9��B\G5���s�iGgc!��bj���-����z�a�M �����I�l�����uP�.Ba=�����
��[_�!����w��o]��>��s��{��RT��-C���*ͼ=�2�~��KM�7��c�|�o�V�����y��@�Ոc���Զ���)#+(�G�G�J��kVz���׌kKi�<s�F��~t�h �^��b�t��+n#��)E�*	�Ēl�ZF�'���&�������h���
j6Z�D)w}d� �G[I����>�V�M���N�A�گ�W�=`{Փ�\��?'�h�3�3�O�#�v	��X���#��I��g�(ȋp8o��R��M�}�FZu8v͢2Dk#_�a�v����LQ$���+�������?J�a��
E\�R+,h8�s�!A��n��	g��%�K��4K�	
��l/+¸��?�E�0[P� 0���<	����&o=�����e�H?�����j)�rQK�U%#�.��\Qu�#�,�U��!w����y��D�{T����a��p�)k	oG*)�)obRF ��A����}e t�,��^����� �e����f�ua�i!��U��j��M� m��0��̴F��?���-�����2c1�\�M]���䉤4��J��f~�O�T�H�tz��L��7f�m?�hE�c����ޗ�_3.S�j�ٺ����GԄE�&�Z	���YG��S#����B��;����&����جV\xpUٺ}����/G mX�-���o�ʫg�c9��릲�>ZQ�!D<d���ߍ�I첀v�c�0Ϩ����dB&'�+~{(@_�I��\�j�E�%C�^
����D��!�c����]��GD�:�0㪀Ȩ����Z}%�J<u1��#�bW�	ht���5Qb�/h��B}Q=�Q�#"ˈ�ա,������mw��w��)���Дg_Њ�f[.stb����O`|����\4�c���"�M�!�1�Yt�U)\�"kfT��'4�X� �<U�X�=ؿ?��짓�R�} a��
�gy�-j+g��S+A�.�T�e����D��y`׵+.��Tcj�\eA!�]U�i�O�S��C{���� =s]���U�-��i��4s�ؽ��ʃ�i���F|ڂ�7L��E(��}z�ݤtk�Ug.5<�'�l�K�S��{��Ǥ���$�����A 쩷�i�\Bo
*���1+R2u���]M;� �]
cʤ����Z�L���&��j,���E=I⥊-@�V�F���Bi���������S]@��ڗ�ΐg��T�����]T��B�G��⹮�h�����[�'�y}Z���ۋ�/%��5�yq��HS�?�0A�\��0)�4Ã�8��S#s�[����7sD�FƗ�	�T�.>_()���Tj���q�����E����t�1I�W�Y��
�	����-�$���`c��3\Wj���t���5�x��c��j���y�����K�:hJZ�!�$&��5��ɚ��� ���yԭJ�C��$�1�ex���[/������N�y��߸x��T��`��Z)&4��$u��Hz�7��T}p�|%�`0��>{Y����`y��
�Й3+y60|�Ǫw�B������e����w�:��`Xlw*U�����e�x�4��]�)�:�CV&�nq����[�33��A���P~�ȭ���iwk��S�>��k#r���	�=��U4]�{�Kn�߭9s9���/A���m' 1eN<RC�v#"y�e1�v2c���l+_fr}`�T�~#G Z���m�ɫ�QB��-�ji(ꍨ�GG>�
`�I�Y��k�b%��uH:�������E��|Y�6
����^��kA��V�'���Z�#2̣æ�֢�Q����_��D9�<E�G7>�ѹ���/�~I�����~��z��o���w����/�T��IJ��hY���Fwt�̻yө>	 }�&�\���1ͱ`���a���ERatK;����!�̻HOFP4w�F����C$3p��P��K������l�l�$1���[f�-�7�m'�����3�	��[3�#���W�����1&�B��T^�§�L���.����B{rL��?��R�ה�ki��9=VK�_R�/��p�s���t>���-"-�4~h�%\�ص8
�@K���A�ĝ�{��,'3������<M�� `q���xR�u��ت�Qx�ܐS���s��RD����K�E]�GYgQ���'�,3��1��^�q{,1A��]C$K0V6���Y�j�j��*�[
�<�j�H+>Z����k�����Dm����}�3>
¼���y��S�wy��G�k������l.x��j`���i����YM#-����kP�X�A���^S�" �������`Թ}Δ�Sn$"�sҩ����q.H�#��-K���@�q��T�z�}\���^�jp��m�J�d���n� Q�[�ڷ|�Wsy�������6O
,6�5+�銞��a����c�LVO�;�k&:���o���q�T�6{�S�����ЂwQ~Bs$��!���u��u�w���!����b��{@�]� T\����2k��i�9����$���ߝ�W�r����O�8�WN��6��F���V8T���7媈�ⰣҬ���h0�q���O������k��	��x|mG�K���5�l@3��}�렎rb�%�\M��c�Epc�+����$Q!�$�����[=�_iH�H�c|0�Q�������Iս�B�`~����(y�腚(�k,�Xf�I:��o-�ļ��y�7'SdбL\=CH-^N�nD.:�X���n�D�>��8=蕇ou�#o������T/�ڧ�>�;q����HO�Z �  g��z7q�	5��6!�u���@|�K9R=_Gc�n\	�/v�F���H��n��9YP�����l��D�h͉��0�5��!@=�ޭ�h�=]-���8N��D��t�.P��1�w���;�5`^��hF5����QMxs�/;ӷ�x��Z�Q��W��߅:������diX�0�}�H�]-!��0�2֩�?\�ª�a������\��Q�Q܊��S�P�$O��Pѐ8Z([�R�N���;�4����}, �7v<�����<sg���U!��4;�h�`A��=ꀣ���;��CT���J/hȡ�Q�(6�x45I�f�b��%Yq֝��
�]6ԩαt�^����e��S���ܪ;�q�1�$��\YE�-P�=�t�syA��腼��Ef���:Y$�*�#B\�f����a���遁�[��Ƅ��s�6�t�E΋�9�8��њ���J�Y�i�!�qmL�Q�74�Sӣ�^�%�y�/���f _�m]8S�?�PE���7��;�;������Ws����l����2���������"��luI'�7�U�R��"{O_�]�G���ݺ=I?`jW[��ˁ�	�����K�\��*�cr�/9��{f�`�#�(�=��w k�cn��\.΂[�9�I��'�l���y���: m�a��$�;�Km��%ڞ�J��X=@\R�g�b21ݝwjͦ}`ُ1�M!��h���xjU�W{� �'�ờ-	w��"/�B7�Te�	�D� �ƣL�|�_��;�o�i�9�)ߓ~�w�cN����uP"\��%z�^}�7M"t���7/��|���m�����$�� �}��g
,P�8��_i��
D*�W雛�[��?�nl𝐌!8�F,�}�����,�2\��:$�E%�e[�s�\��j���Y7(u�WQ�_N�b�����9��v��l�Z=,�Z���m�3�����D�=�Iu,���Stڇ�x��iX%Q��A���Ax	��L��.h݊H2M�I���Q�&WӶS���V9x�n.�̋E
<h,�``�� ��˖z K3!.,̨Ǻ���d2�ל��Mx�^���|w����z̿N�?R��	r3�Fd8�߆%�Z즽QrP��C2k[�!��- b��T6!��c�3%Z׵����m�Me.��:����ݓ-���+�����_z�J҄���0P�@@o����|ƅ��5�B��yq�s�a��`��+_�`9A��d��cm�f��&�~�;�,�D$�h��r^�ނ
V>��йz�&� �Q4�&���Z��O��@Xg�!0eY���w@ϥC*����/�}����@��E�UM�1��Ⱦ�����j�*��Z�JE"���g�ڹ�$�JEng��<^�8�����ʅX���l��>�$!|�;|���JX�[B��KP�N8�)��y&��j�{�28��D$�DE-i�I�j��P����6T�	A*Ƿq<�ӵ)N��]Dl!E��2�˻ڠ���	f�!�pe�Yb~�~n�������ï�-�$y7�o~hLho�Eǥ'.� ����-`s���P������Ā�-���S[�v�78nA�<R(d"�Q��{>�5����.#U���Ř��Js|�FN��k0��U����b��-Y��w�
{�jƼ�ٗܠ���^.sd]�)Q��1KV�<��u���"�o����i�uԱ��dw���Pj��^��j��U�;� �i��!+�,��(��ѫ��Dݞ?=!４��]J�Za���2��[ӵ��E���\�%}��C=-�DI}g�(��bU��I����I竈Gb{n	���1G���T2u�&_�P8�~QwY�h:=�(�Ĺڪ�k���P���_�0-��UзĀ���� ~�!kus�2��k����{���p�/JR�r'.���02��6B7�������ԁﮆ�]�<�EK�?����齻�����*���x�$�����RC �sh�������H=~��QF(|m����F~Iܦ-1�Z~|�qF(EZ+3�$M�b�1(\�D�QbZ$@�Ճ[�nBB��;5�U"���Ol����旅N�}f��XNqwFb�/����/���h�W\E ����T�:��&u�Ճ� �,�M�e�}���k��峎�/����`�W�ZD����m`_C�h�#�� �B^�-���>���Ru�ݜ5��h	\���j�Y1��hB&�R�[�6t�%�q�ܴ�ugm�;A�;����s�`�v^t�{����<%1;�OE�PGΫͣz�%�C�FvPj΀�����ȹ������BF�NX�ҩ����Q�`m�~���(d����{�Ys�wx�u8�����c9G&�߰R���o�s#�Xx�,�7�pOA��q����gX��NJ'�X��(�U�Z}�����H�b٣���2�޴�p����{��J38��z\?�y���oؗ+�.J�?|3�nO�qq��[���k����a}��H;��O߲�I���ԥ��r.��&'I�Jː���s�ju+C ��%V܄������l���	��6�v���>��3{���x�����ܲA!����3��Œ���Z	�V�n��LMH��ȟ89�������Q2���Zi�s�"�|��j��K�����ŉ�'������/�ꬸ�|��;C��f4i������xAM��(i���$L����Yܶ�UӲV��==#�9ݘ���\�`A��u���L!γ�	kqS�.v��*��J�W���%7u�G���XÜ�{��J�+�uL��^�Y:u���L�5�y�8�o��6�j|�S�n�#cDC���F���J�)�/v�?�⑹�?6j+�T�����l}g�?��J�*& �������p ^�0#�LZ �E1{�3#�~�bFb i�^�?)|�4�h$���Ű	J����A�9럾X�������)-��	�p@Yj�f]��ߓ�>�
T"�-6j�2Ԙ�����D�GC�b�},�uMd�o�H|��o^"�t�5f���
�?�R�H��5\�g������V�,���*�^,�:������+��Ɠ�`��x��G��*"S���䀥�Ƽ���#�$�,"��H[k<�_{��G�p�P���dI=� ��R3�r�)�VyZ+�̃§�-�GL���;C�.DUs&�ش�AQ*�93�ZN�'�����fE�������c�>�A��{@����o�@��,�u��������.���j�c��(��+�VV�d���H���kx������ϩ=�*��X�k/0�	���Z������ği��yG����jx��;S�c
�q���J~�HDg�>11��E�D��a+�9��o�<�鍲Q�%r0{6��(����q�-_,Tc�X�_ӓW�a�E��]���A�\`�%X����^����ϧ�JG 3b��3)g?9���X��es����HO|���9\sװ�rT��nȧ�Vf��d�	������|D��W���@�!�����"6w�&��M�t^��Ps�J;����R���Apҏ^��Uj#v�g�FCX!cO��ɢ�O�a��������+]��.;1,e�����2=l��UM���ݣM�?�Ta�D�p>k{7�/=e��7a-lʦJ�tA}�l��[!�B��dԁ0|�ç?��Қ��$��vVW�;�u�EupGj_���*�ś3�C�)4@,�Va`�r�Z$��f9D��'���1���@���;�����G�su{��i�;��[�	ޠy���*)�*q�m��B>��1�C6�fŌA�r�v"�(���&,S//R����ȵ� �EMd���\����9f�w�%^��#&�mwQ7̟0��t� n��s�/rv8��ə��d�j>:	�ū�^s/Yuec�C#�P{�?�r�2�.e�Q"қ��D�ps'���J�;3}0�+p#�����ەc��GW��XbK�aAENx��T��s�f�d�Ԫo��M@u�sVp��L��\���>��r��MY�u��
O�/_��W>>�]�q�%G�R����H�׮���,t0��}��G�e�b� &��c��żШ�m���S�~s@+�qa�����Ym�,g�ՇX�w7�<��a�@�"���y�-����)ۢSq���t��e���BM5r�LZ݊�ϫQ�ьJۯE�=u:l� b5����5������d�����D/�؝��:�}��f:��o[�<�-��,��z��.�6��>3�{z(>*Gҽ���+�ay��RG�a�)6!��Q���W�I��NU���=�Wk'�E��/�H8��