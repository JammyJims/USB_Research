XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����,("�=?��fR+�ϷV�ҩ�*��jr�����>�(4Ch�G�4�_��;�;����w�~7B}e��w:��y�'�9��wcR��0џ4�{�|�E���o1�L\�d�l��kd��5Y��QM*HA�������Z2���ZN�T
��}��@$����COղ��@˰=�q�uK�œ�.XnE�ґ?��h4\�r,W�d����ˁN���!��W4��!#���Kɤ�i���C,X&�����4D.�+�qA��mā$ɉ#�<�g>��!Y�@���Ŧ��,S)+�6������8��O4���}��0��y��u��[l�܅�cie�=����6��8��fng�r��FPa��D����'(�'�
�y~"�-�"V�36�O64ű�����l%v��{���s���B_M�{+�3��y-l�Ya�E����O���v���Ln�C���[Gf�*�h��a�ꎾW.9.S�8M������ׄjx��Ҭ A�Ү^Yip�c7%���1h���z�uo�)��\:�QO���ծ��6*�U^/t�O�_^���8弌�)��'����U��s��)I�D��פ���Ԅ9Qm�����sG��z]PJ�ȱ�b�%�_��+��Q�up�Hk_��R����~jJ@�	Z����5@���j��W�	Bў�@���#4����k#�,��$ P���3���WB�����[<`%���L>]�gՒ
�s{�f}XlxVHYEB    6a38     ea0q`��OJO:�"��%#�K.�;��Jl���Eʃ���O���g�QZ��V,�MJ�}��B�ʲlw��_�N���
�	w���{m�����.y"��&��SG�/[�'4�����p}sAP9h�:� iUV�w���^*� ��-E��~��h`y��� j�m�1������2�5�Ø��T#BDy���-r�l�c�Y�����dg����+	����`���d��w\�rع �#b�W�s*�i��g�&؟j;g�����>��!_����]���M�#�,U�Zbs�����),�O��R����SUs{Esa�[S�E�7�*6���G4��Ńk�4�����8 ݚď�ķ$��;�װ��%��ui��=�&�n:�BRv���]�1����/2����WHx���?nbN	<F����}���zmJ��ziBF�stA��e�%��!R�0��`�_�~�Y��o���n�9dɛJ1��ע�&	�Ev�$�|�R�GIǼҾX�|b���rc�#r�X���R�2E���QF�w���}�
R֣��ߙ"�L�P�}ha�����yX�����Թ�Z&?|�PPU�w��Kx�w ����>}��gg�ֶ�P���������2u�p4�t��&Q��i%��X#������ݵ��V0-�9y;p�;��ߝ��������Iz��k[w�\Y�f��tl��.�}��ބ8�_�K6��1�}!K)��l������?cá��7�MW�����N:T�*����#��%_�w��U{��\�� ����W��A(��*S�}I��Y�h?%�T���� �pT�\�z�g�"��x����D��` �H��[�.���nP��~��A���̓�o%��
�L��PjC�r7�~�s��7	#���Y����{ŅӬ^Y�g�= 
I��wR(xN��FoI�,���&�#�S�_��Jc+0MSCC��|�� �Ǹ���h��ܔ>ƵJ�V
N��
d^��^��[�.e��[�qV���*���Gt��[�Ш^z��z�k0�8�ߺL��s�c�y�/+�Evw��x�gp�r/����zx#jU}\L�}� �TD}0��-�2��q��B:�a��:ۅ��B�`��QM�"SN.UA7P���8��g?J�h�#xyΊ�7�� 
.�Ʊ�9��%<��H�@����ˡ�T �Yc�h���9'z?��y�2�v,�����nG�"�gi�f�h��_A��r�r�;��̶�����waPڿ�XZ�_tm��*p/yђ�m������hi����혾�7�f��0_6�?��4/\��s�p'��J5jE��p��:Ȯ0A�P(��!}9�e�Iؒ�D}_T/'"[alC��D�b�2h���g�Y�0���UH���?)x��N{�oغ<�H���x��6�����o��	B����PòRaZR
AQ;���*.��-�Tl��4�l3><!�����A�H	�T���}��ԟ𸽙���Bvu���!L�?&%�:Ű7�'�j.\�t�ռŐ-�J��@�b2Hh��2oWA%MRjtKB��TLW�_�^���aJ�B�fx	�ĉHY���76��o�rK��1x��N��Ĉ���<[	&�G���7������Ƶz/�/��r��]L���BӉ�rEH��Z5����%�u��$�UC\��rRX�u���l�ш8g��(�{Y�5���-컋�$�A�����ӑ�%�0f1˧�"�8}�g/�KE/I����>�')�4�-d<*����2��۽dR����d5� �3h�Ì1����:�_`�������?�*g/����V�����+:D�d��z����q<������e�K�5�N����a���8U�묙18w:A���pX�!,��,�gH#`��O7�n�2k*�'mG2��6fxe̖����6�pwyE�yLcԋ�T�T���0�JeU��HIю_ ����� �/H*���c�ͷǳ��Ŕ��ˏ�d���f�l[�HZ%�`\��HY�a�%f��	�����}x��fZ<V�|�fQs3��ϼ&m{���t5Ս�1/Э����3Ie���)���s�^��$���=190磈:�okz30�)qC�1��3 �o��� �h;4���5�}�ud���m56�r����]�Y�?�I��=Iô
��S��!��J ���w���?�F�"a[|[B�,ecN써:>��-r��&�B���[���!2�V��}��.N��5n�H�}�������o�=�J�9�=�o�VO%���F�U5�2�KY�	UäBz�s��E6`a���@]HQ�4R3�M?;�d#��f��V�M��%����b�W=�*���G6-,G;�E��Q@��_�wl�>��`:��	3RB�����j�rK�BD���C��d5c�	[>�L�u8;7����^hU�@nf�<�� �s1�y�U�ۍ<�V2d�%��(��ﱥt���Vh����`?+ ��]r��9���Ӣz���S�'$�f�h�VYJ H��=%>̃br�>l��'W�иe^aH)�Q��[��\}]���?֗5#$,t�-���Yd�N'��c]��H~7��.j��_���Y,����n��h��\7u=T�o]K�*1B��)�d���������4�i�������j��r.@S��%�-]��-�s�
��Ϊ�w�V������+p\ nɢ��&��
j?c?����[lBحJ��^�[_�ܷ:4[I�G�s���v/��S���6�%��!���q����y�1���������ُ�ô&�KX)6sƇ��hF{'r~�3%��;�V8�P3������sظ�Y�O$��Y�f��d��~��i������ȋ^��iX��;�U���	��q��;�U�qJ�^�PQ����\�QIYC-�J�V���y^0��2,�&n�+��tO%$��r����r�u�ѱ�W�b|;�����fi�t��I�YRï�۠��\Yfm{ߧ� ����҈O\t�O���0�V���U��v߼��!):�Ǽ�S����OYxG��G�����o������#o) K���>�z�������x��zhJ��o��Y"ڃP�B���x��ײJ�r<��4Ի9{!�t��j�p@v,�J\H2Qm���
do<c�Bt���ۢ9�{O�{,�d3ɫ��ȗU����kӯit;u4�����&j�����.�}�շ������<}��x�z쯑b�:�b=#�+�}��~PY�s$,`ˬmK����}NO�k�-�Sp/���{!�9~EL6���k|��%(�ţ�-zbJ�Of��x�C,��!xjGB�L���2�@�"�l�שӣ����!D7�r�[)N)_W���r���<^W���7�<�8Ek�+V�Eq�T_5��v'���%vu�tK2D ��a,�ц��+t���0�0ٸ�����:�nN���s���n/���X����r�_Hw��;)���L��#�Z6�-4��p�_}ی1%ٺd9&���/�00w�2Hu]�l�������瀣�B����b�]���G��~�Bu�k���L�GA��a'�w;�kY͖���c��