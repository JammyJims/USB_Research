XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����r	��[��dlA6!�4�dMP;G�@�^&�@eRu))��gߝ�G��J	
�^��s��sv�������Գ�N��S�c���u��;/�<��Ma`�����[K�� �=C6|�}�yt�4,��#���D�w��x�T��O���J�k������-P��oIҖ��Җ���A��Gʭ�S��1 ����I�_����o��am�
Ќ�������V�����HG�OQ�\,�Bo0rL�AQ]ds����ֻ:��.�;�*wQu��I�.����7|�Lڵ8Ԃ5Ϥi�����֟��K�#�
�9���M�[/�}J���<H�?$΢^(X�\�-SRf��Aj����3�8�n�Q	>���lf2��l�Ya^gPku.���j>
��;�[�Q#�Q�ߔ5�ˡ ׮�l}���:�J���`��B�����z�H���P�ɴ%񅲉��Y�s��%?K���p���$��h����?L�S���'�]s�e�/��T����qHu���"!�7
Lf�5�n��L��x�b��u}�u�Gi�����h�\-�BV�v}�e�6�]l<����!lm]	Y������]�0d+P��W$�����?�^�@�e�#�?�uN^N�<�?@���"(�f7J�րρ�bkd�B����Y�3����2+t��BOy^���^��䝪W2�۲�*v��A>"]��Ɏ`���D��)Hؐ	��ˣ
PK�O�c������X�N����~���_J���4�z&u��	�XlxVHYEB    fa00    3400+5��Z~4�\����GP�gtӍ9�`�ꔎ�M��Ѝ������0�!
�0�g�"P�s� �*mQ�j�ƚ.��p�Ց��A�ŪZgg�� ��{
<B�On��`;��V�%ҙZ�^.�N05������U�=�F	�0]},5gy�H����4ؓ��"`�*ǣ��JmVq��3}����Qy�!h�!���}� V�Ϙ�F��D��!�%����97_��ME������X��.ڨP���P/��;?O�@^Y+"�欮��9��J�έs�$��p����.1��8�^�����a�d{ˠj��
P$r�k�I�(T�ez��|,�E8�������ힽ�#&��>����lW�;+��T�\_�jR������l�o��z�ҹ�iE��P�zG��;1�u h�l���pxC�+���\wA�t�������@?�U�Q�O"�a���
}A��MF0�ώg�Γ��j��=
��IaPr��m��Ea��&���6'p��B!���""�����h��ћ�
.}�.��N�L�`di\cb&T�2i4Ϛö@6	$|���p�o#�
&�4��[�]�3ꐄ�����n;@� �sW��MdK֩��D 8�k75*C1���|�� �R?~w������3�J���G/X,�~6_(1O>ww�ݲ���MJ$��Ї�Z���׆a��nҶ����Z��\�.�;�~"��0�"}��_���'i��!4�1-���Q�-Ὺ!����l�J�ss�Ϧ۷��d�42��l$�4ܨ�w�� [8��%q0'P�k��a2s�	\�}���m�6��*���Nw�-vu�(mu	 ��'��(ŗ�+;/�;t�Hh(A�ґ����u�w�*o�Y�%1!v�5V\�2���Q �rV}�î%BK�,�;:��+|(�'�ӊ����ZzPRGR*���be8����h;Q��.�8�_ض�i�Q=!,d�,�O��
9���RN"�g+�a���A>P�pd�H�-�
 ����[�r2��Ò53v	�"֬9!�z��iE*���I}Ԇo�,���I4����'	��YI#���2WI�==@P��{��B'X����
��ZI{�x��y��Td��Fs�U�"%�^��5�&n�2��eꥵE!�����BЩj��F�!z�~Lӛ����������Ws��Q{�j�P�rV'��mLVT];�1�q��YyK_��F�ж���.6��T��F�\�RB1�ћ�/�*��߂)�J��# �}����������O5*Q��^�{:v�B�� ��o�)��t%�G�h�� �,Y<� kMk�_L^����q���G�G���+ ̻fF�����>14�ҴS�3Mz���%�\m�|�J�n�h+���l->(L���yy.��!3�3؇4�ߣ`}E�9�_�ztl�a*}޽5�Xa�����%(�EoJa;��oѪ�Y���\��X��_��w�gsx�H47y�m��TA�9?�wAM�g[oЅ����T�
 3޲$K��� @L�W��{H�o�j�E]@W�����5(���o:�����)����|�EW���d�ف�C��n�����l53��3bT���Ԥ�[�Y1Ȟ�Q��'⼺Q�%� ���(�Sׇ�
S�>V��w��e]&Q�>���i�X*3��β\tvx��QG�=����O,�iG���=qSFʉ��ZY�x%Α���T~j�1$`���-I�U-��[Ò��F�[�-|�z��
b^M�H t�1�jRg{ R�g��>�w�(� ~I$�l5u y�oXp5���Kn�:�<�s1N4`͠���Sz�w��ij�F��)19�&3�Pڟ����Ό�۰~,���\��Pp8�t3�03Fވ�U�W}�B61˴ ��|�Φu�4���D�:]ww��Fs�?�q��m)x+o��{��%�$ͰVO�D�H?5�~�5(��&�]����q��ꕊ|�H����j�G��&�FE���O���� {+ᶢ����h&��:�B1�g?���$��ny-�k#cYW�`a`�%\gO��hҁ��.��s�,(F�=�4˟2�`Uw����|�Ǫ
�Z��T9�A$�9<J�v�J�䃜��ݞ�L����͚�XFzz�W:U>�J��\}�$)^�Q��{�?;�KE!��V��}�iṊt"Ba�¨yU�	�N|� ��<����Ɣn��l������9H�@db�������D�:��3�i?@D2��,����ߜ���f�_OLQ$ ����39!5߽d��~�d3�_�i\`+U�%A�	2v�q0f|\��V�X%�zkڕYtH��h,CWƵ�ykI����\�z�o��� �7��)>H�5�0��8�Y��^Z�x�t��dj
�/��(�!R��_W=>��g��I��7�c�v4��uAJ�I ��~�� ����
{a���}]$�|��]����=�V�������T�-�W�2އp����/(S��o� Ap?��_R�Z��(U����(ױ<��:�(R�j�����`r.er?���C�J��8Y��썟�W���r�j�j}?��6���)��Y�RtKRu�D�i?��q�<~$t:QzLK�;��b�)ck�a�;jܤ�>P�)}���W/�W?��$��#��<ǳ`Yl��&1��F7`#m�󳌡ϝ?�4���B����z�)��Fn>�݌TЇ����H�;3��F;O@�m�r��w��e�����$�G(7����\����{��6�7�WI���^�Zh���,V�`�_���vM;�t��&l��"�j~��{�P=���g;�5�v4�Rtޓ�X�5��5�S��4;�f\�@U3�IX5�#��>|��c2j�-�A�'�hT�u�$s:U�����*����̼��ԇ�	#�,lK�0��޵A���'<��?Ї4zz�>O�`�� ��s�~Z�[Æ��a��dI[�;������������]�I=���)`���`����ғ�6�s��;���O]��{�9s<���$�S?@��<����qP9H�G��ȵV�R.�x˰�d�?���0k9g7z�7���P��g�Ƴ�=1^[e��#� lWre�)!�dm i!/0��� ����<��+>�L>k	��j_�`:T��Sn���2�n>�Of����=�ڛ�a���%�%�D_CV��&�.Z�t���z�̽�=AD����_C��zѨG�;���x����#��
�*�ݜkHe�z�h8b1�����\�iB�d�B��S�9)�S�_��N4E�og%F��.�'ƾ*����@��\Ɯ2�$SڑwgK���I�����'�\{ ������a|<
K�\��w�4�'�q�T�Nw�6��3Qkc�ٺ|��0���_��
��Pi�D��:����?h������dy�}��Z��	�`��A��܇���Ο-_y
���t��"�)?����C��kD��fo�P�R�V�`��j���J����������ע7Be�X�3� �cY;�@�]	[�	�'Δ�m������>ڑ��l�`�MťXB[nC���趃�:9��#�:����⁯
ʾ�+T<bwr�x�W���yER� ��f��fWJ"Q��y;��$ο�~<t]<�ӳ�;|3c�l��/�k�U(fQ�Qn;[}�p��&�/����V��;y������ܛ��W��_��^2�2a}�{4-z3�4�/��SJUi�t{Q�����k�Fa��	��Qg_�a��]5���b%QwO й�&��׎ >^07��Ϡg������iv p��-����\`p/*S�pz�;0��blSrSAc����MNJ��Z~��-i����goh2/�iY�L�ۃ�g������d�1����͋,2/���͓�����<s�{��(��]��=��FG(
�7P߼��=�Q�8�S}U��F���zۀ��pV�}���\��*V.*C�~{�:[𸏥(�K 
�Kz�!�m<E8��4e,P��:0�ſ0Q�ǮÃ��x
$L�ȋQQ~F^�^.��v��ɑş��-v�X���˒RM����6	�&�M����uq	뙄"2�V�?�+>g��Fh��ˀ���AѢ[y[�ܙ�gKH�)��k��a q�zl�+7.FT�]t��1�܆w	�p_ͅ�B��\F�n�M���bC:D�����z��6�1��bE-H{wu�*JE{n�fN8��?�������*uO����k��Lgt���9�N	�H�0/ț�[w��X��Kʈ�O�A�U6�/+�	H�p�]�H�Ǔh���s���g���hSV����k���.�ܸ�H`�8�}��Q�T�~�*5��S��R����yO`�+T���5��I�`��QM�8�B8WS��L�nΏ�zϢE�����k ����=TS��?�n��1{S� �o�S�*j��īP_	���Z��C>�����WJ���]�\p������y몐~�O��SR�;������C�8�M�>�6� 7�GO�6�2A�&��Z�2�5D�t6������ՙ�>܈�O(BH_���m	o>z��MY7o��w�A����|(���ۆ�PNwU���_�@��0'ɮXR�B�H��68�K>),��
�MJ�޺�sf\p�N�Ʀ��K��!�w�h�b�Nz��d��ҹ4��+f��*��ę��f�5�������M+x�nrL��`��}ϸ���*'�jӂ���ʬԥ�i=�7ce�ر�݇��#��,��6�	�7��)�������F�9����b���1��h���E�&��xy��Xׯ�R8Pq`6dwG*v�x�cj���"X�T�j<� �OτX6���	����ͼ��M� ^�[c۾���4�Cr&@ IF��l[����j�^T^�5v�z����8�6�Q;�+"���ǻsV���(V�aP0���Tޡ�IMݩ��,�we@���WRf
��5-ρޚ���TN�&:���e�HT���ܡ��KJ���Or{)㠧.��Ti�٨����;-�E��OA�?+�f���l�ƸV�Ј=^Z�H�*r;��wK=��X����13z�0+�W�̨�y���WFK���#���Bt�\�D������
�)� �3������cu�.,ұ	��nG��3!T��2�h�)V�|�0�7�U,�VǼ���o�dq&��LC�P�55�b�nX�m|�S��^v�cA%ka`]���h���ɧ��«(-K� ����B}=��݋��&F��_��u"{KY2��{Mo=#i�\���V�l/���>�ڈE�Р'�D����+��:Bv��D�f�	i$]S�d4W<\enL�w�Q+e�6�,�~�[)D�[_�Q��:04�>���\��l|�R���%�\�'S%���@�4��غ{�k]غ~Է3��K�����'��ڦM�ܲ�av&,EfCϚ��w�B���b�]�ٔje�;F ٫�٣~����1�T��䑭#�B�?��ɬ�d�<���L��P8j�Λ9�s��V��:n�6�1zM'�������EZ~�G�l9w���ǿ����û��J����}���G�L����:��4H0�����s��)e��<����D�*�8��#��	�t	��Lʯ�8X�o���O��K�ضW�[]��Fm^�u��@{���}� �:��p�������u�c�����J@����-V1r�޻oZ���S1��8/�k%��č:X������&W&�0P���Ƀo�M\x-Y9O}��{{Ӯ��`AdN3}
�8:�Ƶ��V�"����%.9���J����nY��j�?�������jڰ>\�)"��kcwaE�>�`}�">���	�'( B/��p�ܫV��7�f@f̶�f��{�����Ngw՗�Y3\\1�8������O���46$b�!-B=���`3����I�,�LU~{��@F��P����OT��PR_����k�ኪ+�Us��d�� �N� ��{��5%ӁS���!���Sɥ�o1�Q�����ҧ\˵��#&�,sz���E�����Dɠ�hDʤTZ����T�`��>��%7d�E��Fk*ǰ����^��[:�g'M��Z	�Ӓ9�y��k�O���
M]�q]�-E�BORN1?������˷=>P�|E��H&riĞ=�=�v���]�,����������!ۉ�O[�#	��b��43I��p�ճ�R1ӊ�S���h����.K���/{�h����o���L>�C+����P�� �!�PD�2��ږ�0dd;��h�-:�8�tS���3V[<�&�E��#$����)�Ⱦ��ī?/=��N�W�C�w�+bx�6�U��9��<XȺ�����W"M��1���Kr���o�Z)��
{2�=�XDo��ACH3�0n\/�#Y(�+GfϘ@���B�	ۿKD:��������w�ٍȃ�#�rؤ��E6���q
�����3�����Q�d7�'�6�E�i��7:>"��s�`��J;8�� d��Ǵ�Ø���bS�Z�0�?�8�OÐ,'e�=ӄ�#
,*�g�e���Ϝ����P ��9%?܅!�}~I=T�^ў���aH���RY�̃��:�T����Q�/��O�A}O��Sk\�������5����{�BdT|�)5��=h�Bl��8��$i�%J�06T0�ŞO��\��+P��7:��&p�T�r͂��PH��\3Mi��M6������|!yy�c�Ct�1�垀�uK��{����m��Þ�6�M�gહ)�������'��&��8���Vh�])��. ��KD��1|�+�;U�' ͎Gfȷ��x2�������е`#�p}�|�9׭����zfi	�*\�������T����H0��w��vs�vH���*d��K�Ք	�.�b��j2�3@D�
�*k�?漸�EW�Q����v���2����O��>���t��+YW��N{K tb�*V��ao��_r
i��p;1��3L*�֤8��.ah�����@���m��.�ϋu����	�
Õk����[X��
r1����M�����L#8�t���;^ �V߄ArH�u�<ꙇr�g��,x�i��Yn��W������̌��ēq����P�2��|*%�~f��v�G�Xufk��6�&{b���ϝ-a�N�����;z�2^{sA�z���]Ϧ�kG������A�ß��K+��H��N%�I�+�%m������+�	����UKTS�[�$Vw�[��	�y9��i�1�?�&��"l�فW���[j/��t�|��/�å�;��Ό�o��Θы_EV{i�M���EȰ�m	4U������Lݔ��Y�-}尰��Q	��	��I
A�&,�N�p3��~����mL\L�uT�pGp,{@DhD�X��g���vt�����5շ}��%g �op���.���w�_3=O��PΌaY	W��v�}5eݽ���,�b�!�,��w^�(o1�O�������G�<���y=��5�#anr�#�})�|��"��'�T^�>�d_Po�.�m���2��~t��x�~�-՟�O���@�dR��ē��t�Lf��"4s�g-�ZG�C����'�k;�Eԓ`%9����->���e�/W4��f�]��ɒ�|ؿ�J�wY $�9I1?q�?&w)7�&+!/�6n[	�e��0���^�J�rI6��)�����{-����ɒuMg�b� a;h�}'� �nB=7�/ps��H�I';�J.w�B�iEp'ԓ~�`x��aT}v�`�l�p�'���p�^���ٽ��*���y]	ߚ��%Tj������̈xs$�YV,���x��b*ٰ��PZ5����	�����U���矷���1\���Dv�����3R�*{��RE�GN3����9tL��+Ž����!�n���JBi�n~��s��W�ʗ2��n㭿�] M<To9'?R�PAH��W�l��f<A��J����g���J���iԧ�6,xp��m�p�W7�32� �T��`����������ӄ1�=�	��S�1<Rx��3۫/+������]d���@"������)�Z�KJW�h�D��L�֮d�X;@�G"����%8z��'�~m�29A9$�7���K1�V58Hr�(ĂS���MY��6DQ�F_3�6�;""���{�-�d��}��Ǫ����"�q���S��2��i7�{��^eOf(�8����U�+��#��K��&xt�l."��1q�J���TB��g�Tc���(q*�/�*�i�N��d&en�׾\ǰ�7�BU�0F���؂Go�o7�X�ڎck���[͠�8���)](-�Y�%�+&b�(P��C��֌���k���Z�]�;4���/�?G����M��/%[���q�WNs�{�'�Ƿ}��4tk�)���ev���I
�	���!�;LŎ�����Z�r�lH��="X�G�s�+�"2(mq}�~n5��Q�];�׌�M��4���Ww�D��Z�mc��%�HT�< ��!ਯTM�u��?��ȇǡ�|�Z�ؕ�#l�����x+�%U�����N��?�6�K��Q8�� �1��sb83яm�'i�ܒ�a��1��qU+��袄Y��e�=L|�HD�d!f�.%�u���MD~����x2'�qPf�"�W�M��ҋ�A�=n�����A��$�����;Ɗ�Qu{q)l�ݎ9�kgk���6b �8���@VU=;#��YP��Q��5k�L�e�T�;�U�(�&��W8�#�.�>W&}4�,���+������W��!��R�����3����E���j����S,���jU�U���x��C5��@�4$eS��eʕ<���[05��15pY:�< �$����(D���t��Z�9�,�uӐN�0n�"U�q�=,F�}�9�>�xV_g]�R\!��b���=��Dà�b�BsTz
\�e�1��'A|�o��M�]E�� z���"���{��3Q�c�Ƥ	$���&�h�t�Y��O���?��2�5�f�(gh[%dK{�<L��
zN�T�_	�U�:�R����Ĭh��q�Ɯ�B(�^�&A']�E����=�Ff� d?;w�jg�����_��8�H�.F��t�k�~�����{��[q�i{n�S�k���D#�������/v�VCQ�z�� 䠪��޿�f�V��2�:�< ޣ�#̀����%���2����%��@D�A�m�
�T�g��L]���[c͊ԝg�Og���bSHP�V�w�ir{C�������ރ��c�,������C5�m�*:'��3�f7� rE#�"&K鳏�S.�I�w��K�w;h��4!��l�}<�Z���C�L.�hUxA!��Z	�f�ؙ���VJA�64��1b�ݦ~/�zώb��%��.:��a���ܞ��W,��/��J���X� �S�>�]\�XX�E�W��1��ul����:%��=�>����. �������Q��]�y�w��z�[����o��5�07��<�W���#)��� 3<]kc8�%,��1Sx2���^Hи�����M [�@�nid�P�	ǡ ���F���K(=�L�۷�vBj��ni#�3f�_���	Q
�l\�g��Sዹ4�J��Oda�[jL��t5f�������Iq�hk���~�����XV)%���L;����V�(ѫ���?T���������=��a�F����Lv�
J_�������Nk�o�"5||j9�������K�]�F�F��ʆ��].�,�70�PY��s#�@V�Rn<B����6�Il�ϐm��ԡ�������j�����R)S�}�Iض\��ɿ��� T?�5��g�5��x����Ut�R�����Z�ַ����Mc��.����#�Z�FaIC�&\~T����E�g�]u-��G(��o4a##�D|_�Ī�6e?�0�����k:����/��K7���1ue���{����]� �TU��A�� WUí��\FL,L�H{�B��>!�(��a��[�<��纜>�D"�m���Dsb�BM0�+�	�O�7�=}6�1򘀈�>q�^L!t��Δ��6��?盰��4�}Y�����U�cD]� ��:'@��fq,ʖ$��,�%�!�����""hW��R�0C�A���'_t�sm��Q�c���,�{�+W�箪g`&<��,>�=&�mōL��4���'|�;��A��IR�e�N�sD�ƨ�k�9@�T�����j���u!ͼ)6��&��8�P���0��kwJ�&=h����A�� ~�2`�l�za�_�o��p_�꫁���CD�D�����v@�QL�H��鿙���q�K=���Ff��)���'UcN(o�a�V�������iTI���^�h�P��I�ĺ��b����JE<��p%C���j]^���p�FbQ� +�a0>�Lv�����}�1�����ڗD��38O��pd�t�E��M��) �B�4Ɛ&��H�;��ƀ��[�f�S�E�b�#��r���������{9bD�q�b�!�D1�o�s�7�O��[}�Օ��G��)�f��S�+q&�����qv,&2tM`[���|�����}� Hnq��.�}�9?��Gl��1����?���j;���5�>��cf��~9ќ������c@�h��0���n�kz0萗+��=�֯,\U?"���à�/���w��{=g�H6ȵ�Wv������ꌘ�X.�X��Lg�Ȱ�K2ȵ����C�Q���j�����k��� צ�J�{'��S��7��;�����h8|_[��O\�>�霋E(]|��<[�c���IV5���4���P�WF7�x��6��8bAȭ��s��LP6J ^8h�G@�_lPGd���-oY�1�b+�CH�C|	��5f�;�ꦪW�W�����G����4u.+ �(�%�W6���mRq.�ʱ�l@����`�G�ʈ��g�ć|S�����$�?j������{�����?2����G��m��ϖS �Ρ�o��i�aX�Ǘϱ`�I��V48��^=/�:���Uh��1)�_��W+s?������RDֿ������������CB��U�{#�ߜ�:�	�j�2c�/�|aa���g"��MD$]����n��;��J~#f���~ڽ�@h�a=P=/[��3v5Ij蔍D�F<<��NI>�\JP���*!��4�)i-tBv%KP���ht}���#z\z��	�����!`�Bj='yѲ2?}�hݺ�I�yTJ�����#�[}N�ˊ�y�rx4&�2`��C��>/�c=�C�x5镸j���J�J
�0�W���; ��$!yj��4fA�a@�+&����P�rݦ�y�k���[EX3w{�џK��g�Ò<��M��fL�c�7�����È��ń��/yشq��8�8�&�	@1���N{��B�/��^}D�*h{R������p<W�q�S)�L��{�@�CAc�	���S%[H+���79������Ϥk�)�4�u�E�̍�)6�S��NR��ԍBi-u�DT6��qbL���z�����z���D��qt�_4��Z!-�������[`��#L�A0��`^)� ���\�rؔ�N�Q���R�K���x�B7��w�W1N\>@�>����'(��č�R�k��c�O�5�w��w�e\���RLp�rΕ��n�,���}�|��<����rj����ߏ�-�zXr�����+bz\�l�Wo`��UB�h<�.���ؽ�d%���פ�Q+�&�Ms��:��f1�j�ػ�<;��Ϝ˽�����$�u�>R^h�>G��B3c�*� :�r��?�4����z'��kh�%c�B+R#j��U�����ڂ�ex��U�.�<Ȃ>��z<&N/�w��������	Ґ��Y\��R���́F#q+x��:�3*�����Ff�z�s�MOp�������N�:�����Э��K����{p6�tH�$)����s���*僴w��\��E����WX�@[XJ�7�^)��Ɉ�o,F��:�ܬ)u��u=�6�=�&IS�$"�E�,��[�L!i�H��:nH�`����ЇSf^3�B��y�)b��(C��m�4]K��X�iѴ�����4(�~��+��r�Gg�����y�3a��M���+Y���m�x��D2���ЈZ��x�1��d��a��;�3Td�o�����X��tcq�!���;��8+φ�>�~	���"��ګJg/.�ι��Ǉ
[0�*�~>}X��~��덎����,O����;��;����l��6�\�I&ߙb�K�|&��>S�	bP6�T\�H�R|��p�rC��v}���〕ȁ� �|R)w����>#��a��7!f�E`���=J1�>��v��s��$��?�x������y�|����{e�]����Nlv���[���.'�-��u;�!]��CElQ��l�@zj�U�Q��c�ɂlz��X���O�1Xo��)/`�z&/?�MiϨR��}A,��"��^��RC����d��.�܈	��=�M��sD�A_�t�IO���,|hQF��M��?r0����Ȯ�2 �0��? 7-��[,�}���
�`,��
��-�Smdv�-�i$Mo��nrN�a�ŀ��|�D�� gG3�>�U�G���U����"h���%����k���Hl�+�#��q��8���I�?��͝��(
��(�1Lq�U��Of��Ħ@j�yJ�a wJ߮ZVW�f0I�WxK����#��V���$L��}x�"����k�
���@��և�Q�+5_|_T���R�P1z3�s��b�ۇE��TI�s@])M�+�!�s�x�,���]������8�§w������D�V]��TG�w�V���Q���Z?��)n���od�z��R�V��>a�ϗȈ�:��� .�S�ġ#s`�-��O�T\�V�`����y�<YXlxVHYEB    fa00    3480t��rX�:�ʕ�&�<Y��.)It�ž�N,WЎ�:e��V۸ξ���tҔ�C:-V(K�52��p��@p�As����0}�sU��s��
��Jrs�y�&eA@֎�G�2hB�<��;K`F}h���!=3N�qK@Q}�g>��m��M���k�5�S�q�6��h�#��]a=r�3�!P]J����g(9_��E LZ�QΡ ���<*-�N7�;u�����%"�F��Ke�Ak}�K��O����'�hR�E��Q�6��Z���=�d���1��鎆� =�5Mb��د�[���%�T�_�-8�������ዹ7����6��@qT{TY�^ �@���O>ǜ��wh�h �,P��t�0�?�S���N��k�Iq�
w}%�@�����|^4��-�� L%��(��x�k��B#�k5�4�eV�MGKfˢԣ���;�ր�\d��tGZ4�D$��(����;Ѽ�gWXR��ȏp*�膗M�_:�`���P�ӌVi�Qu8ھ��d\WA�f�%��9l����6q�&�7�)ww W��:!_2+����Û�-k�ʛ �\є��f�o�q���~��Q�WK�4��B�(�
֏�l���z-6�C�Y$Ib �"/ Q�w�cy�2�^��F�u��]}T>��A}�&96B�RZ�[�<ja�_!��p!�*�b��_YX�R)h��BmU�~�eB���E��嬜��+��j�r��B�%��%S�ӆ?��n���C�,���9�^/
����H���<%�C
�f�t{��-��8V��l��8~g�a,����0�D��W�����%w���}�޽6��dj�7>mu�|o �+W�����0��!ǋ�7��=��~�Ĵ�� @)�M25 �δ>h6�Ǳ��7Yc�S�,�~��u9�	'5��y=3[kge׀�w��K�$e��Y��MW[é�����W胄6K������ig�Ƹk��
�5)�M/�e I"�YZH��t�	�˄o���`��N����`�^���4��5�&˼��U�j谴�PWo������7���'�X��^W�&tRo�e,�Z�]�5|����{�4X�/Z�mY�^�M�l���3�UqEH�Ͷ=L�&A1����[��(��}n:x��W.��7����,�FS��L��H�e�{����=��7�}��)N±���85(1�񟞜>�;�!ҽ\/�e&E����:ǀ�G[�����/�_"_���<���4��H y
=�D�)�^�r�̴�3�j�����+!���2d����9�8���[&�"z ����^|%�z/�x�7�ؓ�h?�5�MDg��v1���m�3<W�2�u���++��{����u�ELH!r��'&��.�-���������T��㛣�n/�x(�!��&^[���?�R'��ڃ��?�s� ؾ:(�b��̅�;7�c��At��$*�S������&���R�8��?pc3��40����R-�i�j�h׮�[3�/[���jDk����f�I���5*6�PF����x4_�qMf���|Eܢ����ԕ���5��&; ���飔�!����P���etW�Y!��u�(-��Īn\�T� k~��7J��GR*� ��ѐ3*��UѬpW-�aT���ۗ�.��9ٷ
�	���nu��=�)��7F�i��Z�59F7�)��i�,"��
o�7���l�H�3�k܏�L��4��*ԭFY���a���G5R�+q6��uO9�W��"ݖ���sZ��?O�P�qjF�Fɺ8�ܕ<��'�!P�9JC��ɼ�74�^l�˲{`���h�
�;��v�CN>���\��
@���i�o�Wv4A�%��N����ԆYA����`�5�v�L�d���ɒJ쩊��7��
}G%E���d�_���& Ţޮ158qW<~z���1�B����亵Ǎ��G��dO�\�\�6 �����V<^�^k��j��6;���#|�`(�m!\q�C�g�.�*x&�x\$K���?��?�ED	��4?���e�T���>.���D4/2<��l3�w,�9���SZ�����Y�����q���'��Ys�HS~�[����=�P�@7���+��nm�� ��<�l*�i�����$K��"�O^K�%Y�,��l�sVc"�th�0�`]X":�T��>���2
������G�c�'oՇ���Fgݟ�֨�*l;�y���Ϳ�����ɵ|鏇(�қeg�n�F 7�enA��H�-l}}�t"�26[���H����$f*���
�͐(P���ST�����E�M�1V"����L�~�l��Q:q��hdҡU�����D6#{,�6 8x^�O�|=�p^+,�G�o�w���X+���NNzh6p%}������d��$��L�4���v�eޮm��B8xLs�?HI��8�;K��*HV�I����@*��N1�[�l:f��F�H�4N��K�* $�2)X�������b��7�`sX_a�2��\�F]>	M�X�r�8j�ǂ�M�4�\ҿ���G�Y�Z؎N�L�������b��#��Pٸ�Ϟѹ�i[ۻ����QKH*H���F���tn��B(�y~�Q=���S���-��C\Gp�⇕Zt88y^j*ȇ�K�ODO��b�����&�f&�* �7y�Lp��&Ȃu�_c�WR��}Q(t2�C/
�)��W�C�R���e��z9G��ǝ��!�a����
�;�����j-�>�4��B\������Ki�G��j?76�������3��u�_�<��Z��O�â8(_�r���9-+���9�ߒ�%��O@l;���I���\���Y�S*}'*kԀ�Z3�v8�Hf�C,�å�í�i�@��)�'F,���}�9�.Y)�)�3ugd�_<C����g�����ޚ��Y���9�[���T�5_ث9�RϠױh�r<���"ÊG�e�|b]q����Ag_��9�;/���?d���)B���������"r�g��yE�pDW�ǰOS��:'�t0�AC�Gl)�X���rO�pI#�]�x���r-\��4t�q�6��L}J���r�R�z����afY�nT����ش$@+��QQ:�  �R���ٍZ7o�_����򉢀�T�>>[�\���XA��m�&;�)˶�(j��˽.t±:C*��خ(��l\DQ(���3Zkӓi�G��a�76w� ����;��A �D��lRZ��Wm�0�T0��<t]�R�눍U��9z�zަ�Ѱ��vh�5�	c����y)�����LE��I<��o���PM?iBw3t��[(�����)���R��%��l�HN������ì�Z!��;?M
�}�)m���ݗ�x�̣0�B�0 ������2@&ˀ��t2۟�qqK��"�����|G��c�DݢY��)�������y��Ό�;�(IV,�+�w�ϓ�
�a݉��DPH;bT�w���۹�в�� ���K3~0F�ށ�`%>�̫4U�m5���P����3[��q�T_ ��K|�2�4V��fĢ�6Dϑ�co=���";��	�[3"C��=�Z���I�seT1�T�(�l��S,ɝ^d�9�1m\�g��&���E}6��\���tr�wY��h;q����;�~n5 �P�:[i'`�e?\�B���<��7�n��{�����,��Z�%��X)	��[��Ph���S����(�vT��y��/-G<�Lps������)�$OF��+OhwC߫�~�?aڈ^��',
E�1�%
��V��Î�z�����,�=�%^s��0����N�<R��4;١fU��<�f�j+li|��.�f�7wq1:���x)-�nZ��K3�������t�x܉pt��+o��ÄD����2�D����>8��<�]W��2���_��m�K[�g�\�YD�15Hy�0��If�NUp�����/�:�d���wV�x:�;!T�E}�t@0���ln6�4.��_c�yF�	(���6���ܥ>�	��p7�z�OK�|�5h��+��"�i�b���Y��.*�ؕ?���U{�L4�8�dp��'-�'Q-Iּ���+R�\���ܨ�XJxX�D�^��>��e#����t��ީ�t`�lZ���\�%������*�ɩ]o��h�<=��� �]�B��dv<_�WD�cEP�x��̢ȱ3@�	V�I�t�dM�e%�/�q9[�D]Nk�m^�H'���k\V2��Q��d��6�~�jh$ݥ�!<�}��I_�\i�jj��]��C�~���@�Ƌ]�/�1r���x�0��Z�2����Sp���bs��I����_7҅�2�ºoLm�{�6��|�@>N{�ٙ�r���B��U��(�g8����A����G�o��h�c^-j��z�L7�>_�9��3�vhΩ��A�+�.��T7�O�*o�c�;�iWk�KBh�,�ֳ�a�g��xv\'TPf�.�q�!���9���~.W�ġ�є����s�A���ё4��O�e?�웁���g��v���Q�n��qp��[TQ6�+������1ln�(T�vZ@��m%Cm��J!��V�.7�M?����O��9U��9���jf(]b���q�(��+��N�r���2�h�p�
u�dM�c��Q�4�VQ\��4s��� ��Nl/D���.���Ж>x��J5�bq,8�5�;�'�9�By5a0
��4_:�'�c�{u���մ��kÅ=��g= ���j�+�*_Bp�a˟�8���y����d�5���G�_J�(HlZU�|g�J�(��/E)d�Ī������-��e��Ur�k��^� <��1�[B�X�-R��GҀ`�;�B��9e�}�����R���i8���l��J3D�o���XZ*"Zj-��b�Z��kR�!��3:��S��Aw��^t�e�� �$w,()��I��؝�e�&z�c/�y�U	�V��$%��U��*u����J)��#�p����4�u���ߏ'i� 07=�n�o�~bHa���٪�(���Ι����f�ӵ�7������IU�.�]�g��C.KS���T{���Z�����vq�g~b �+[�vf8Up�8V�ě���yK`x�s�u��d"'��'�-N��N��	���^���2���Ӱ0W_���Z��@��T���I��Bge�u����o�&��3+!-5[&��5�?��KU��d.����j7�s�m/l��E�����#��`�᱀���=>�{=�0��V`�7�&j9Fy}(��#�㶋trF)�+�� ��0ˆ]��kk�'�_�Tl��Uʈ=L=X�>���攐��;q�\[�)����I� ]0]����g_���+��m�*j��L7�8	cn����ΞI��o&����f/¯��ͣ�*��K� ��\��F�O֔K��H�!�2\sg�ڼRZ%D�#�} ����ɇ�P�!�M���S�#Tլ(^����@ -4{�������ڶDjV&�>��zq-[�߲�7������.Ws��99�Q$����f�y�>�Y��*އT���}��3���z��{���(�����e�c6k.y�'�(�op��t"
�;ɓ74LU�q��&)]G���eq�����3�l���4|�њs�
'�$E�ݍ��#�Y��Ԯ��W�2-%_�\3&{ϘL��v�Y(��̢�`�~�K�'���*������Egc���<��(_�݃��)"��:���,dg\<�t�y�<��n2By���f|$B4X$[M9��uk�]�0��f(�� �}5Y�ro2�����;P���*_���=t���)�q�t�x���UP] �7T�QR~�Tz+0��N��8���i �!�r���VЉE̓ƪ�m%9;B�m{%��Rz?q���ZoL4:�>�w��OuF}pn��ς͟���r��d4ى�1�F�C��R�� �gk�E�E�4ÛYe	�B��s����8�I���������@f��qíPR���p���%�C>��_�𗡚6���Z��4�?-��E�鱚%w�Z�RH7wG�w8(x�\�u���0�_@{���R�a�f}�	�����Cs����������a�G�g�w��6���5(5�a��`�|���C���T:{�g�P���������A�O����8���%���B�=��C,ʿ@���<	P���~�Q �B�*5�~�+����~�9�p��A����X!�M,�m��Jl���M�=��P"ͦ(�N �A��b�����Ja#h�F����rm������=�����I\��YU�~IϚ1M�dl+�2Vn��Ūח�,�E�b�U"��UW.�g��B�|�lD h�̈́���t*��IXD�5��P����[� �A�<��]����8z��D��`�;�����X�Ni��T��U��{���?E��~b��K���d�e��j���j�g :k�z�:��[û�xӎ���U��<频�V�35"�p~b�$=%�z���[H3���
I�_�S>�P�^���U��$iE�Ǖ��[���u5
s[�+��ƺ���a����q=!m����'�f�D�z�h>�Զx�Ķs/�z�ђA|�h���}�ȳ�__�-���5ܬ
i�|���3pzb����v[�v"�����q���\VG�(�}E�4��\�UX<�ꖋ�ض���P�-AX��hA���~��@�s�>g{�m1�/]	��Hâ@�v�S��M%G:��w~f�A�+��2�A�M��K�����U_Q2_e��`D> όV���s0���yV��o�ԗ��	ʨ@�]�o���@oU�V�qm��N"�m���#���#�2���M�!�+�P"�t"}���6AOhl$�8����sW2����Q�)R�] � ��2i���,�7#�Ȥ&������,���Q�ۇ���uq3���J���s�1���rY���CCM�#�f�d��g��8��?��1��i%���AO�M��c���I�F�F�K!39�gS�ŀT�V�m������G�3s�V#Yx���g.J�Į��ί	�^�r�� 0@�w[�B�c�5ټW�&A��``��՛�����P5>�O�����ڻ�_Ӟ��'gm#{��7_q���gݝ�Z9�v��mz�*���cBE��>7��!2���]d ;u�� �}�:L�p� 2�k�#�PY����EcO��T��~�`6f��'4�~`��X����~��¼h���U(��t�%L/���+tOo"�b��Y(�6��yJ��tl���Хa�#�ϕ��%aFыYa�2c��������l�G|i��3���]L�]rKՅ�(
=�B0@�k�����tqP?���U��|4)�v�2��o- �tF(B���EfP��c/y��h�����T�m*xd'�բ�	{}��@A�����1-�?M9��L�����������x�G��ơ\"/�S��"yhCT�����2_���KZDu,����	���P3h�lG,#�&Կ�Jk�z��?')�6�JL�qۆp�"ĩ��{�#MoCe�\f���d� <���7='#�>?t!/�:~��P6�L|�����CQ��G#d��2£��OP0�Sr:6���? c�ܬ�{Ҽ[o�����n���@"K� �]JC3���ION�q�>��`$zf�^����>��|"��5ɃܳF��-]�\����:����*RU�C�iQǝ������`\C�c�d�E)�4T�V���b#7�u�\u%QN�
����3�|c�Q|
�.�apț�?�m�7Y���~��u��>x���ip�D��O"BQ�xɎz|��ڳ÷�}[�s�8�٬+�4����DM|z�����Gӱ�a[�xr�� �ǁ�a��s�M��z z7����Vt���?Ax��Qu��HRƹ�΄�P<��z����jS�ٕnN�����PN��}�a���9pnk�P�n:F���@iefr�z'�+,䘘�c����vU�������	F�T�B�x,�9S
�f���Bެ��Ӯ�>�R�����H�p�D�9��4���a�"�W�� ���[MRw�@�K��	JZ@ӵr���(�éP�����H�ɷ��P/x���u�˞��=\�v�e�#��n�V��H�&݀(&�׍Fߤ��hM�z-�4�}J:�&��A��s7J�r��_���o_�sl��T�N[�-�хi��y�����.��U+�# w
���/|���+�tV��Ƹt��w�<�d|��6�;LB�u�Ėǳ�ێU��O�1gեt�e���M���	��A��õ���T�����Z��3;?ź��7Н6!�ֳ_	��d��;�N�Wrf��_#s3C�S�-�"j�lf�L���m�ew��n��k3ĠUwn�n`Q�MaE��қY_+��/�zu�;��.a񘬆���:��1<�q��1���X F�u���l߻J��V�\���t/l��q��:%e�^nj.���z�� 9�S
x����s�����5�50^R��PI�r���2A��L��'-��T�8�|�pQ���z�Uu�jz��gA���0���~u�op�� %�98�<ϻA�5[�/땾/��g�?����j���C�[]r!�����h%��j�ʜ�w��u
f5�^�P�q��"����}Hp�?L��D�8!�ﵩ���(5�����^��Sse@������80%Ȣm"�G�Gq�I���X��q����'�KԴ77�GU])��״�9�goB	g-�N��o�-�B�-p`�O��ޞ�`�
�5Bg�5�����b��d�z+���Y_$8VkZw|z��N�?L))ץ���4= -����R�}}`".�\�a�VQ�ŔʎS�`�7��D�'5v}��koT��qMޚ�Z�
dXmCü3*]�5����٦�~ �
����U�>P:��T1(�F�Lޘ^V�̞/��nlTS��e�8�w�����+p},�؎��C
����&Ξx?@F�9����f詽���C�4�g�Էe�c�(~-�$�6�bQ��~��T>��-�
1���F]�?�=�cf����C)]><Am$8�R�W������hGQX��o���B��';�	����Jr�$�Z9y�䆳,"��/FR�Ը��#�D�[+zg�T'��c�l�LN{�]��Evv��;����� ~ �%�GP8������}\6?Ĵ��i�&)��#�d&A�/B�.���W)�|N��p��_�:\���6>�\=~�N�$��9�0s��"�X�ǋ�|a���,s�d%�&��jy�@K�M�.F�ehİ'��v6f�0:�>Y:��#��ò��"�UIK��$�ͣdB�,�r�|m2��e�p��(�5�bS^\�6��r��k8�g|�-F\KR����\9���ѭ��m�:��C�-�>�N�6b�)=%-_��`+ݼ�t[�ʉ���L݃X��2��� F<j�Ll��b�_u�"�����s��]X3�]�i���	�W$I�79s�c��0�zԞ�"�d�Ng�us#�Y�����)Z~�4! �iqB�+4o*85d��AP�̡�/��0o���v��ά�j�߀��� ;��庐]R�C��N��73}_'��6\���͜�-��p��	�RP-.8C�|�)L҇����s��k��S�Zٻ�Dԥ8r��.C����c���\�vue����33J$����k!	���ty����Ay/��lh�<+��URH+�����:9v%bW]8k%��z"4�0�&O%�����qyta�D�n���)�:�桟{،Gr�G!�[樹��DH�B!ǆ�.�bb�&;z\�!��y�n	�(8#\A���Uf^H�g˞k��}~y�om�bݨ��o���N�Z��v�5�H@�eW����?vv�o��E��s����]���F�8�q�3E������{�%JDM�bPהp(��g�G�����V�6�j�Ms4A~���f����݄�pj���(Z���ގ�8�l�d�Q�3Y;��ъ�ٖ���Gt��t!rۗH�sV����MN�g���T%�!���O�ܑ�m&�ǈ�ʘ����W����j��a�ћ7}��+�޽>%��'�jt4Q$�PV�k��x+�0aˮ�Cx���������]�]#O��s^��><�ޏ�/��g�����r�(�B�9�F�>�&�{1\~P�s�
Y��.���8�m[���q�p���'��;fj�h��v/I�
��@��'>�θ�i���'���ܳ�a�w�:�4W���Y�/
��N�^��L��m���ɭ�$/��#$�<�bS{4�8��oF�BR;�a�b���ٞ^'M�]���꧞�j��T�/�E�ա�a��?���{QZ�I3�1\A$1��it�hĶ,���g%���}�Q��K.f��[ %n ����]k若�/�S^��+�/��J���
O����}qAݠ�^�ĥL���q�x�5�@����&~kme���;% 1p�����T؞�?]1`
��YTd1�F�v�4�h��:��`�+��B}@̔?�"lRx�d4�G{�-���0�N���34�_�jhs6��7��W@QI�Bx�!��ۏM�\�]c'է1���� ޻��W~"�bG;���J�t��Y5�m���P铃��u�mf5)ѹ������G�/��Ў����m~�F����ܚ2��t��4f�n��^A ����������C��.A�`�'LuT@
�	��<~[��L"&�>+�jˏ?-ߴ
I% _����g�s��)���p�����O	Î�f/%~��Xn����V1Ȣc�L9Ǝr��g���t�m�8/L}���^���0�����%�Z<�h^���{ ���Ąv�%�⛶��i�O�.$k��ZЖ7�� "m0W��1�R���Q	��P�`�h�g���lL`E���94�;�[���؝���Y��Z���������^#�L�����.X59�Ҥ��p��&��f�7G�Y����x�T��xՇw�t�(@�+��+$a��á;�@����rR�~��[C>�D����ʷ�q������R�����!�.>�3��χd8��uRkHGcm���������|�aZ!�`e"����U����W�n9�g����'�}�x�.�))�Te��ˤxdI�؎1c8�N�bzQ\����]f[+�
}jzp�{���kg1���q��-6��R�����!�`B�خ2�h�6�d3��I߻Fn8�.cT���߀(Y�)�Q(b,#�)3��H(� �*�}WY����b�4/]Q�W��
���J�V���f�"/�9f�������m�M�k��)UO<�;���j���u1��^����^×[v.���u�]¥�_,��"!����R3s�iͧ��es8���i�[(��	��)څf.9�T�������{����i9~u��但����T��1y����o{$��4	�s����`Z.�,@���?��@��CHØ뻌;�v�E,�vl"\�<��Q�L#abք�R�q��	 C��%��T�gGkc,�q�Թ �ů�PcC�B�~pM�CӀgĮ�D6	�vU�g#Ӵ�zO)�u�m7Zu���-�_��p7���u�x(D�{}L�t�Չ�vL*���ܪsB6�@�����%~#���=�b�HRݟb(g:����`��l�s'��K�U��<����w4�Kj�#v-O����&���'%�f�e�NGk�er�X;�,���&)�</7.��Y;��8 �킵N1��/�a&q��ۋ�D崳&�ӼT����4#?�3�L���n��EWVnu��>Y5*�rݨ�����wP�~����bo����u����+�������U�HW� �>�y��ô�/�J��Qo��b/R҈	�ъ:�����})���㫑=#�����߯�^C�����!:[v���r#�(��cCs���-tF�����;�a�r�G���v��܍/��c�����|��4���k�>�+(o<�,�؏8�&(ōr��=�VB���|��8*�by�uC+���"�2�m-�S,L�o�pڢ5{t��☝��Z|!j.޲���hI���/�5%ȑ�fN��|3ORHξ��Ͳ$��M3������~�������A*6VݗI���ڏl	mD�g[&cp���ڧ�Ƶ߅���+KJ�[���x�������U�nF&/ў��O7c�s�Ko{�4'�x�����q��ދ5� kx,2��������3��z���p �ߺg�c+9���0���a!3=�z��6�T
��蟞+�'~��� �bA��N��$�1��T��l��;��
&%��&)K�g�J���G��D�e��#*�(8���jR��|���cj[��õ�ӭ����&����D^{���*4�I�%E�2�˗��^qP�����}��-QQ��<���W�v	Ѵ�&����&pǌW�{�t���6s�85���RA~I��ɉ~U�IҐ=�w_�5E�p��x��T�k����V:{�N{���w��v
ׯ�,�oJϰZ���=���pɶF��y����x�?L�?z�aK#����ch���s��-���Ï��$��T�i�PI�uq�/�f����Lۥˋ��S�p�@�~a6ӡ[���&g�/�H��ؼ����NT�W�����)��c׌��y߲�FBkS���z~D�����/�C�S��H��~��5����.�����/�&LOb��S�|dL���ŘW��$j�H�jJ�c�2@���M��?�4�뎅�-D2O�یê��e<�A���B�17>ZD�ʭ��@E��`�@b%\�3��I��g��|���_Z11���v��"b&C�H�UiD^�|� �����t��������.y5�j��I�^3�p��y�9��M~��k��$�z��Q�r�T)�He��$�u�&!�*q�Ŭ��xҍc��B�{���M%�<���o<H��t����~����k�� �aR+3cfA2���c�O��󺨮�%�Ķ+,��g4�n�1��޺�;a�nHXlxVHYEB    5980    13005�y0*����b���p��]����,,gxa��)���$F���P�ϙ
G����↗
�u�4"�~V>R`�!o^�s wո6/A:���F7xSۨ�'f�2&-�2t�d��[�P&L�_մ('�	��^��M��D�����5�G�S-�Ҷ��6�~f=il��>/���]�$}���B��D����H�<n�d���ځ������Ͷ��,R"T�	U����LOWm'Y��~ ��In�vܸ�q��Y��m�үT�yWd�j ���9c~u�K���f.�.�d���k\�6��dݨ �P�Ҝ%�^޳r%1m�L�(�g��������g��/�P�(��% ;1Լ�5�W���!�M[���QN hm��sځ�^�;+�u�|�fw�A�苮�ωB\�����ݸ�P�AJEZ&8�B5�L���c�(omJ}�&ܜ��3q~c\/T�Y��R��ۖKH�� �-e�GN ��u$���6�6�p`��Za������Fa�\O�_|I�$���/*�u~!�c�	�P잀i����u�f��C�X�O���8c{N��z����.ۥ��ǷI����1!M+�>W���K��̱U�~�ۓ�	'	�
vNq>A�ζY/ڞ���!Rܬ�g�Mxs|Cs�tP!MS�F���5�$����i} ��-�]l\���>	��M\N�]"�"�*SH£���2HM��ÝdV�&�z���!�-/!Z�GұQ[n{��x@/��x()7�$%S9���Tl��(s���4Ԕ��U�}�D+�.�_��`�2�2��ݹ��!���N�ɊH���g̀B��\��,��K���J�@$�ū��G���^:�T�87�B�x4�'*��5�Y�J	ƼYx}��;�~���!�o-!���ޥ;	�!���U��\��d�,�Npܦe:Hmzz�>��X�(���^�7��K�	�TM��lO<Sa�Z"-Wa����'uP��X	�G,��+*k��O��{��O�e�n����/�F����q�����,�L��{ɵ�̗��{A��m�P2�j���pX#������'��zh$��ur�J����p�.׫��V&:R5�nL]�D������'�b5�zeHN��j�i��߈�����݆C���u
'}�V_��gz�j�qH tW�91{�P�r�^��ע���~���u	Z{m��i}/��ǦO���C^	O�'�
TE8LE�ғK6�'$�X'1c��WA\${�Jʰ��#�S�L����@=���rU��[��qh���v�z}&�|�ZG��aQ�}�����X/�A6��j�`��fϓ�U*КZR�;��QRtp���0z�ݑ-�u極9���-�Õ�81#�� 3�#5�]{\t���=5&��{��ط�[[5�) IҒ�I��s��?p�+����Ʊ��.�MY��[=�k�ݮ���H�aÑ�m|��8����L��K<0�Eı��'�'qZ&ڹ؃�8Ĳ�K�#<J�zx�I���&;cn?)8*��_�s%p�|G��pJ����M��*w,��:�t���Cyy�� a���xs���|��0oی�5��۸����X��_ �b��Z[)w�9��լ4���.�Gݧals�S-d���Û�P�T�{
����%�Ǹ@��\�9&��������Lf�r*6�Ô��b���c�3�a��4���ۙ%nB��D�{�Nt&50F��m��Jې�)�JV��?u�������(q#�62z���U� �8!��61�2T��'��{)��2P��s�!y!��xs��Œ�b�*���?ق�A��9�B��~<T������1$!�-[E	X�''YQ�e,4鷮���3WK���;�Rd@��XGV{;�.��+�V$C�KU�݊�6%�X�Q����u|�2�[a]�g~~&�%����T�wT�c���߃4�Z��{�-Oq��cR�K7sc����g���4�=�h
�0̃��E����^e!1?߶>fWa᳂kT�1���/f�PW�Noc�!`Xi��d�vz�TD{Ц� ��r3���F���5�KᔏzK瘅Q�7���>U�k�$��Ĕ�����
�K�یk%#~�����:B��m\�֍�Æ>-���:'��A�ҝ��5��'��w7
ҵ(�z��N����I[ʠ�:�Ԏ���x1�&))��c�,$i7EY_)�)M@��n��7f�������7���_s���Ԟ+�Cb�^��zu�� �/�\�6�4��͓b�)��U�y�ӑ�T��p��ȉo\��[�Qr���4A�@�Ӈ5_��N���b�U{^l��,�Hc�ܸ���,�3!g�@�u����`rT� ��*í�f���=���"��B�T|{�����fZ�bR@c���-y�r�q	����m��C%��� P%���g�\_��o0Y�-	>���,���pK��%��Ug��.	X����łM��_%&�Ͳ����~�+������E_��鉇7��cgn�ĹD�[F��K����H/�S�^�#�s�&�������uw��s�j����H��O���{U�aE��>���ΧjC0�v���,X(�v�Ӷ������I�����hG}���a6Ĺ�ƥn��J&�ƓĸhdR���>q�F4/���C��6Gm⿔�@����}A[?�`���_�*��:S������<�͜/a�I���.����Z}*�K.Lʇ3�l�wY��T��D_���O�J��6�[���3��&��o�/�7���ͥ7ѳ_��:jy	�qZ[�#�l�y��kh�	�.os@4��#~�����}}��]3tM�r�#p�t��0��#�[2�!�(�L��j��������[ ƣ�;�)�'Mc<�ӥ�8s2�W���=*�'9�>�O��$"�`H\�d�.%l>��{����~O)ث.˟y$�Nj۴��O�p��X,̓׋�0w�T�ooe����(��͊���c�'���X/d:z����8��y���b��ht��	6!z �_b-I��B�h� ��va��«m,���f�r�i&�к�XC�+Yq`�-N�L��RY�K��Ϗ�g�:�����v���;l:J$;(l�v����i|tq�����[祉�K�Ag��ϲ�s�%�K�Dsᔗzc�p�tFⱹf.w5Ū!Z�z�~}{�`��� �yd3:&���r-9�z@D4��{S0���E���>''���	����U@2�ݾ�௾�;Pƅ��H��W��.P�f�b�u^2A*�D ���W�R*��-�� �K~���y�ej��>�_�5�m�f$��P�A��A��؞+5:�pIm�k�$gl��?D�f��_��N�$"v�F
���i7����͂���=C����P��gU�n�p�`a��J�bEq�Ȏ���<�$L֮[asS�N��[�i�ƍ���h��+Ƶ�kf��X�j�>CЦ�
6ɽ�g�����$=n��*�fX�h����3���* 4��\w�n����Go�_����Z���<�.�ʤ������w�%��T�>���<i����1�����[ ��.߃��4L˗�����Ăp��5_�mB)�⩽z��/�$ҍe�@Q�/�ɒ���niu�s3�懏>����S^M�b�tωd���Iu���4B�X5}j�L&�Ι'7T���֒���w�8rI���=x�>�^MB�����{�j|;�*cc�
Z4�4��Q�q��_�mЬ��A�~�5�������5��GC#��/CPռQ����5������Ѫ�9���!��������2����n�幪`��PM�,�j���2yv��Ϣ���k�V6�(�Ԙa���m��!CU�џ٨7�=jh7�|�F���$W��K�3�D�x+S�w�0��\ݏ���O�{m9�f�"$bk�X�w���p��A�y�[·�-�v��\�}��"?h��nT/:�F" ><��`��(U��cv�_��ؽ��5��-}"*�;�|ݜ� �-B���<A� �:�� U�����|&{�(S�����a� �;�$,���E[>� ��9�����=��P,�t�!�(
�1#lX3��$g�i=�u��o)f��yd���������<TV���E�� fJ��̗���{�_;D�&�y��,���c]K�s�p*wJo��e|�%s�@�2}	�Ԥ��pm���3�;� �z]�U�3+i�;�̏f�@R��v=�Qb
��k��¸���L}�������B�l�I�n6v[�L��x��R�c�]$$'�#<�g�Crg;��Gm�n��>�P���b�H-��P�HPj�J�Yy�h�t<Ż$�!�I�L�JL�d��"��C�'�pf��7��:��Ӎ?MB	la��@����0��:��6����gM��f���a]qi)���̴���xQ���4�����3�j��3v���^��h�"�=(+��)�J��I:#`���iQK%��wK����0,�%��L �❅|.�wP�J�pY���*�V_���DAt1�<Xo��3��+&��̤��v�ɰ�Q�!U�N�F�0sVa��_�S�B�nP
�B��F���_	42�b���"<�=�M#ж`�P��\�2��r7J��u���=OAS������M�q-%���=n�m��y��0	G�������d�Q�f�Q$ij��f�+t�9ݰ~Kǳ�A�R���9���H�)�M������!��s�����T����ί�
