XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ƿ&)u��f\���0#v<�!pߩ�E�z#�KB{}{@���V.:��n��E˄X#69U!��F �+j��[����:�G{  ����	���ìփp�â��Q�ykݘ�$�boYn=��藱Is�C[Z����Id��?P��N�O�:�ӟB��_�O�� �
�u�I��i����`�^g	@��2�a�B[���ko��+�a�v�i鏪0�(���L�<��J�
7�#�C��r�+B�����՘!V�XP�V��v���y��ȕ��y�4��Ou!�@Z��r&�m]4�voEtb�I��0O�V�^������?T	fov=���K~�W�)���7/�9i�)$W���.͛
9���	�s�o�Տ:�$�A�z�Q��.5]������1}]w��E������k�ި�סJD�0��w�*����Í�^�W!�#>wESi0�"��^-ק��>�x^�L�ݏ�X�gS&����O�HT\�F���������]��ڶ}�@m�����Ӊό��c<�:���;9����\-����JEiǻ��7�T~2�o�Jgڙ&�����I4� pǖ�@#"�WCW�W<��B���E�O�E�?XL|�dg\[kQh;���ՙ��U������C}���*��Z8wM��M��:j=�vȇ�H��qj�Сۍ�vYj�KQA�bXz�9So4˗D�
F�B	���~��Q@ߘ��}�%��$I��ggI.*bWT�Eeg��^�XlxVHYEB    fa00    26d0j|�J�>���k���c�"�p^E7��1�
ye�}��-M.�S��l-���z�n��d̖��H7n��aơ���\�ķ(��a[oGe�}ӡ�%�8O���������Q�[�&E�U��į
g
���.���/�*��Zg�Ō�Y�BՄq6�<x1;��;>�>㕤����������+#����De�	O�@o5m�>���_!i�5j��7�q)��0/�K@E}ثR\e��F����U���IT7{o�����W_�*k�v�Q��\�+/w{*1�a��w|��,pf�@�r�!�u�B*�嬰b�
#i�A&#��^���E��������(2D�bԵ
z���J���)�5�e�yDR��3�5���G�tD���<^�H�Q�D�1���ʝ�ǂ�Q8ٿ��}m���~�!����pcc�dR���lˮ"��!Y�w�C�i�A�Ƶp\�<�����y�U�J"�����>͋�{ǟ�w���a���(ۿ�˩��'�������G�AT'4�W����q��m���AP�K�7 ��eB�W�ۣG�U��[�úfq�L}��@Z�ҳ���2�� eK��f�F�*9>!���0���^c{8����_ǯ"�O�Vy	FOd�=���yN)�BR�ȸ�Q�1vq��xE��	�@U#]�*��ݓl��=e0��W��{��9�-�=w��ˈ�ex��T�릘�~�T{v���W�P���I6�4�#p�فZ����r�E0]*�bXxҿ��a Q�S���a*���E!���|Q�Gc$�-��/����K�y�o�
�h�yjl���3�����)��N)��c?���,�j��+O���%t��:�d�ݢ�SΚ�12����=�ؤ�v���@W�@�_���5��:�����Z�
h�|̣����q�|♈�X��c.����}5-�ۻ��Eh��(۩�q#(��妭��h���w�h�����u�ғ��l,�����3�K�p)RΠ�r狀��*�W@z']J@O� �.N�b7BZ��k����>�6��,"$���J� �7��|dY�b�]o�-�h��{s�#)-9P�'%r���)/�2'��8�(����\(4OԚ�����ڒ9�g�r�vL䂪29���uf�����Q1��9n�k/(NW�='>����P.B"OZN���I|�>�����ڈ�� ����D��i�aJ����I�f�������r�2�$"R��?������b�%JUA����)������JB�L�����,�&�E�\=F�.�KLC*�t�(;#��9��i�M��d� ɺz�ۄ�����&H��=\&c�)�!B��έ��#-�5�c�e�T+�	�P]S'o�Uy),��j�x#N�܊P`w��
�;�&K�$eE4�5��� -���i:�XM�oF�׆��0���V��v��X��7��R�檅?�}���hu�0�-ZUQr㤚lE���oT�ѝ(`QyEj��'Bd�SP��Md�Y�6��}�/g�(�v���c���8\ !�V�8'���.�da�I�1�(��[�ͻ� �X�ҮYb�CF��[B>�D�p�W�����$��a��E���N��Zb���I1�����)@Us��V0
w\��ra�}2���Q��7,�g��-�	���M[/��(z|��,4�P��'���P��~�?q�|���9F1���o���Fphg�t�	\���'A,~c�ZC��*U��G-!���s�Q�jdބr>čd=�&z��g8������vLuL�$�Jq��v�Lj�ܪ�a��}=Fg��L$cA��Vq>��T�FL� ;�?��&F�~�<e�
y`	|q:^�h!�25�9��������6W�8�7>a�	c�^)����%4�H.�[<�ܼ�3�X�V��e�p�5k�|b'�)�>I�y#�k��Ut�{sw4Y{zM�!��z?
Խ���\���]~����9`)�Z�.{�a��MJJ�Hc�F��{,	g.��F��!�*�{�ح_����Y}\�Bl�ɜ?��`�_�>�Qĵtr�k�_��P�5�I%9^1 Q�DN��~N{o�=!|xS�g��;+���ip�}}�ַ�pw���uS,��R��s��h
>��E���]�2E,���r'B	���k�[���^��cN�4�dC'Hd��Tdr�sK$��غ:�'u^�MG�kGc�}Ut2w�;T�/��p�_�/�ȩ�����6���o[�%hۏ[i�����:��9K3�/-��j��4�y��y1�m.�8��K F�\���Y���;"�I���	,kZ"�׹������4��5��{�⥐��B+syvKc��m��G-=�Wm^��URNuQ���	P�0�?@g��Pe��p�u�4�Q�ϧ
Xvr\�l�jq�R3N�����q�Ͻ���f�ᎆ$���}�_�1�+�R���c��Pd�$���Q#
"��o%�5�U1��F��FTZ��*��vyf��$��f�$#k�\�0t�E��Bq�,X��CWZ�g���Wg�2R'[wq'&L�ޓa�B#>����:����+VM�,:�(5GH_�7ΜP�`W�"�N<��f(nQq�Fy���NF��K�SE����o�L�3���.����-�˶��ӧ��bρ�O�L�*Ɂ"[�ˣ�w������.Ѣ�o�l��>[�y��&�Bu&���k�8�+�M�|�^ LFR����Lȗ�'�>�:~�6����H0����{l5�~<��{/����RR@�Ln�ٸ��)��2`�������N6�V����P�|Ǵ�S�ǭ�ر�"�E�wE�2̛4����[���z�E:�~�|�|��W�r�&���u��S�x+�*�
1	�Z�k�����f����3n%��L{`	��MmL�(�
^iR��?Ć [Śe\S�e��p��v�p���@�|�m���S����y��r��( ���*tT�	��^����I+L��ƖO`��A�t��4{�ϕ����!IΡ�)�v`�,ܠ��F���8��L.�h;K���o�)���#�6D�t0%�|F�}��qS&�8,d*���?"�P�8g�t) !UQwY�N��V�J�v	�H+:��R���$Ҥ��#��;2 ~])����k�v��������DM"�k��.���Sș(�_03G,�/.�1C��*���7�2�+03�`�K��j��T���G+�Fj'��s���G�a �L�g����^�q�����}ל��[����!݋H�xtZ"yg�����tE#�(dbi��6�uA{j���ۥ�"v����!��S���z"��A��T� U�'�I�a4/�	0�(���!J��6w�w��[f�ǘ0� ���t��aQ��]�5P��� ��+���Z)n��#����X���o^kbQ�gU��I�j=�H�O/��r�P��AjDa!.o���9j&� ��vm٪шqn��[��@�k��%_#p��Lr����=<�Cv?��t�'�dj�h����D
$z� �"���Z��D�G$[�Z�B��K�T�S+y41u��	Q�D��؞��X�.� ��o�<��]�x��W?\r	�s�#�A��q��)�7����1o�@|����j�:g=M�j����b�)^�Ȏvsiξ����h&L.q��*$z5���Fã�_���<��m�(C�_D��T~�g�8U�偉�]tx�\Tփ�}��.�ܲ�cc9�W�Q��.7i����#l<�=[��֚�a��W/G�&]7�9�%,�k
�x�`�?>��Tc|J.8����|���#�7��y$����OH��l���v�26�QwN%�"�,HrV4��
\(���)>H6���eQ�sy`�_�k�md^�$�b8G�z`�Fq����s�Aୂ>��s�"+Ӕ棄_�VT� �������;�d&+��TC����Ԛz���y��?ߣ��E����A?���y��x�d
8o� � �P���C#޸(�n:�"��ɱ3\6�7��Bơ�K���~�c]<�K�1n`�W�����J�d�k|߬K�ȯ��E�'���$ɤ�s�O#&��4=+� H],���r����A�r��saF�����(tkZ��.��0�����KܖΓB�(5�<N�vfc���A4;R|pY%ꥆ�*�C�ǜM�\n�::css����&`L��4� �D�İ�3"΋�����)�A����_-����XS�7"j��Y|b��L�[��>3��`KzFM*��(��HPz���3�}�������2���i̩�q����&
]�^���&9�fJ�#SY�a���#�w:ʡ�<I��4˗<���p��W��<N��ZY��͓���xMSJ����h����ڥ�z�Y�����I��)�0�9
u,�P:1nF����T�P���pG���6"f�`�q�aS���o��!���GM
���F�����<��g���ډmhi�*b6k���9b]C�`�[���3zy�M����,�C�s�쓪����v�H�tYhQ��Re��W:bvF��I�M�XkN;�yy���a�J��q�{���6���HAv6A�뷫��&�VnJg%�����Q䙆������Ռ���(�&�I)�(	����)�*fӂI!.�u!y8u%X�H���{g������N�� hTOVC��@������$}��f5���}���v"�_ƣ��fP�%<:�	>+�#�H�Cw�ʫ�\PG��_w�c�PH;�P�a]�h�WD���b��X$�_O������7m�B�Ҡ���.����~zR6�G�߶/BIm�K����q��E�C��	v���H��ys<�ch��.��R��l�O��6�ǳ��f����A���7�{�CS�9
ul`Ã��dA�(����7բ����G��-��]�VP/��'#� (Sm�h����9��+�� �0�Q�c.LLL]B�+;S�h�R;e��$��!9o��	ќo|t�`Gv6����O]1B�|6KX<]�Z�h�b	��i�	*�T��%J�Y��l�e5��d�,��2�W޺��J!UXj-׆�����8�l���n�o�N��tzR�:����#^�
�t�v��%�37Y1�b�2j��Wę�l��( �E�ԁ_���@��+��ħOU�x��Q�l��gg7�Hi�.~�Mͥ���N�'~4-�im2=������dU�&O�j�\�]��XH*�_�QpniX᢫%��bԍ�a���N'���/�_`�<�AZ�0Ϸ�ﭕ�0)ve�_i��8|;ȩ�ttrɻ����\��n�Jv�*ʀ�On$��J	�����syG�!#�?�XBA
[�����T�1�����%����L#��1X�}15A��y��K���ӹ�������
R�.,������a��K=��@�L9I��4]����߂���L���\�Jl��z]?�Ek@BFmo#�;�ٔ0dU�w�P�H�o���$L���(� ���c���,�e�2�gv���R�酘U|�g<�B����Wg�l��ٕ{��ӿ�!�:���s��Qp�(�O��쉒'��@��QF�����6O�\�h#3J�4��NUo+�n��ew�Pz�@5�l^�~�}��� sR����צ��ԸaM�i��z�[�FblƠʍ�C���6z������	b� ρX�@%�B|�@���]�]�Bؤf�/���]�=�&^�r�a<��K@iD�IBX��:ٙb.Փ�q`oǉCa��0�I]��� HjaoȎ�1=�@:	�^y����y���Fa�l���4;fh��M�ٕ�'v>8q���sLQ��3[d���� 0-�d��]
=��j���)�p����H�z���b3���f��-6dޮ�[�H�*�L�ʄ D���B'!v��]�l�w���l;�߾�Y��,�!���������>����� |����� �ڟ ܌����(�oD@m3���[%�� � �8�	tz���>G�ܼc�@GkÏp��Z��HH�g�����8�Yz���"st-�\d����f�1�Z4%�6���`[�n�/I�96��d���������z1q�����z��[ylG���k]�n�4�ջ�0�;~+,�Yk!s��Hl1}fW�Uo�mԦK��^�]Xq7�rt���O�U�J�2ۓ��Gs'��#viW�f��40�<�;M�k43������ٟvٮ��{yHT���u%�_$o挋.�]�\�֧tz�|���4���e��[��HnS[�wr�>����5������6v1z�Ǟov
�ixr�G����F笖�V�Q-,�o$��-E�n=M�v�[��S�f�������94�j��ڛ�J��Ҽ�F�}
��o�ܞڻb�$x�R�o�i�i�\I��U^�OΠ�\甸�N��Ԑ6l2g�{c6��t��ݹ:�j�t����hQX~��0�����k�"j���e�+�\uY��Z]�R��aw���]���z�\ԽY$TٲK�4�$���z�Y�L����h	�f�Ѵޜ���8��- r�Q�(u�`c���H���Ԕ�G�Ot���L���T/�<(Q$$���ľ����ub�n�G
��6�!\X��p	�z�:Ʀe��>�ۂ��θ�l� XR�ʸj���8d�(F+���F�gf�e����ӱIy�0��1���T@�C0V��Raآu�?�f�?�Sy��'�=ѧ�5�>}��WL��v�2�����;����� o���3܅w�m�R �ߘw4���s@�p���9�O�3���O���jT�%�}21���k��
�_��W3��>��Q`�ʚ�w���&��:H鸴��ȃ�F՛�s��R�
V��!b�_����ф��g�������>d9s]!-$�� ���d��={�i�8����^��iE4�/�-��,�������&����L�����6�L�1	���q�z.#?E5m�N8���Ǩ%�]��k���u�xa��}�����-$<k~��U�3{!���P!%B�類��`3�|Rx��W����©T.��XI���;���p�zP�V!-b��\�Z�hm���` ���D"9�I�a)]��#Ѧ�\|���7�Q}�︷�3�[gŘ}��H���B������<Fe���e"�|u[U���R"=|����)��ர#6/9[s�R�# 6��q�84D��ϋ���l��!��>���Φ�2�h4@I�s_I��.N�P�eI/Te��R̳-�/.{� R��3M,�z�H�L�vY��
IT� ����X!�H��� u&�[0E����uQ+$�ҹ�$�<�x~*�'��gF�&nP���i�D-����������8��7��%�[����,�Y8U0f$���'Y��?�]A�����?��ZUչU��;2��&uK�1O�����r���C��%K�Hj�I�kd9�F��!���%į�L�9�I �&-���D?vY��Iє4�+E�~4��G�k�������d/IV�k����vÑxӃ������P������H[��H�W��Q�v��w{=��"dXl�H�x>��&�p��׏��t�~��VäSB"�4(M�f28�ӂn0��-z�똄*�%��X�r�lF��A�L(]��+h[=vY(Kj�-O!�)3D�^�d��M�]埖Iqu��v�g�^6J3�a �������;�;�X,G�]�:Hs�>N �ؚ�3fvvwbʃ��WY��R�ۑ�zp׎��	f�m��ߖϼ;l��x�T�ׂ��?l�~�-	P�$��=�0"R�=4�^<��r�Q�L��aL�[<P%�Q��
��09B�"�IX�k�����v��o�p�.�Bђ���%݈l>�	HH�c��Y�v��[�a<ҧF�,	,��6H�^��q�n�ަw�nK�xɿ�%���t�v ��Sq��rp#(j�d�E<]	U��=\��BL��J��T,j��N{�s�fϙ/�����9��&��޾P�y�B��,G�"(��-��I[wC�9g�R���}�ߔ�0t5��b�'� u�������ޅ�8�8�B�פe1�)�|�����V�]�!�uU?�������-��&üS��*�3��$�_��ԿD!^\6���p�Y|�	ABhx�m�M�?>v�6���ݟ����8�@~ �[
�]ؾ8G|4��2oJ
��>)Ɨ��bL�Ĕ2���f�9����[�ѐ�{0/qq@y��./ƮA�MK��f$����Z|	���[�Q��3�1����8�&�K;?rT��\=�E`��.`B��Ԕ:��Q�����r�k%ndʽ
?'M�6�~Mrm��?��������ΩF��Q�/�n4��ջb178����{��р�cy�o���k���'�CG+���[���������\W�hL�F�N�˘��+g�T
�|�	�9����j'.�9�����Jm��aH$I�\� _��|Ņ�⒃�{���ͮn46�����m'Nc*z��y �Yvפ�������O}�Ǘ�VE�����u�Ш�Ng7��c��e�&S�)�=�Up���PR;�cb�O��f���DU�$z��������Q���-j�5�F�q}+�%	R֔�2���u-JQ��̶����z����h���א:T"h�����9����(����u�{�|��t�آ�<M��W<����J�a�,E%�jJ~�Ɵ�&yZ����t��l3=�wxPh�(V��M�כ�/��i�-q���r����� �ݑ�B4fK^����Ef��A�ʏ	�a��|[aC,Kj�������'`�z��!uĘ�'�5Ӊw�!��t�4��D�G�.��iE��,Oswu�l�҉G��q��>���q_?��܃7x����Ϙ���$��[+��"-��WFx���RĲ��`2����@2���+m�?�{�N=Yq��"��Ӣ4����;`�ٶ�E܊�,��~3�SYw|3�l�����.���
pl�s��8�Dw}��B��\�dǘ7�V�}��Mpmh�CS�K ���N��k��6��H/�3`�
�m�����7��;v��q�b+�V�B�=��l�v_��)X�T�[�'d�쳳�
�S�͒�Zt<W4D0��@�bo�z�;��]��Y�����C�"G����p�R#����˫�	�m�u8]����=�(�V�Qd���0��|"W�ə��1��\ި�#��Cd��6�R�`�g����%�����t����<S�6�~w�")4��[�.}�}�l#sC{/~�%u�� ��S��8�6���N��i*��M�ɤ옊c�5ņb9OsU��߬<�Q��Rߦ8�U����6��>y� ����&���^�!{��S��^N\h�x05Ӿ3����5�R�x%;b����_�!L�\7�������R�	�V�X��fy۫�ڍ^#`��>�с�|3��������5��<����Jը��}�P*nb�û��#�Z:��Y��Dk&_cΓ(~�Cd�A4�IP+��dQ����j�����ԯ߆�QR�_۴�![㉑��V����9�4:�U&�|Q�'#��r���g��C>t������H�0}��d��)���}�D1d!6£�>�I*�ݒ��<��6`�,�
�W��������0(>�p7 X�ʞ@����_�Ν��Tn�k�1G���XlxVHYEB    fa00    1050�#*�����>n+rG%E�A�!!�h��J!�L]��~���=�����;�N*[��(�儙Tb��b@�}V���)�5w��z�Ɨ>�G���=)��PTX�,c�揄���|�	}�#��'��؊h�?^&�+��@���z	%n�~����%�5iN�q���7M�]{�C��{�}�q�B:AmER����*L����.�C�-�wĳ����;,��+S���Xr� jugyl�~nˈ�At�&�c�Nx��5��֋4��(�I���!e��穀���&Ґ��+*#&�uXW�s(o��l�=��rLf`jZ�WR��]@�*uq>������Ol�	
�y$��9�y6���,����?H`��|3A�ik��c0I��J��C��6+X����F���^��1�m��%T.����!Q�&���U�=����\N�o!������p%vc�0�˅��S��	W�!W�
�VTɘ ''T��5��:Z�5F�"���j��;&�/3dן�,
��O�O�eD�aV���-�?��j.���D+(����a��ZaA����T��Ov�:@kN ԋ̊` �����U�m��s�kR*8��߻���bhL�4�B���X�)��������0ٴ�P)O�d��Jn6�ݑ�Ct\�S��4��jzj�x��x8���[�+�wo������7�q�����V�#�=e�O]�������su֖�=���u~{�`.<���_�Ae��NRa�䀬J|f�l��+Q2�=U���&�_�m3�G]�/��3߮�fl�S���`8��
>�����(k��Z���81��Sq�3��>�/��Y�CHm������噛�O��-ς��K}�ޥʡ�f�$q$8�'4�Sˡ�-_��YJ��y�]���5�ϬV�K���]�ǿf� ��%4hq�.����
g�U�ȣ}^j@����M�k�E��GX+n�c���%h���e�Y�C"UҗO�x�ZUN����g�����v�Џj��4�ʕ+���!_�>�֋�g�j?���
�^���y�z ��hA�%��n�V�
�����:l��5�%��8>ǓD��v�W��n8�x^a�!ζi=�D��*E��",��D�{{M��.&('17�6�&RNNfJ��;�n��T�P�"��̈́ޡO�0Y&X(���J?GEL�¨P-=�~�fhN,�AĖ���-
�$�__�Lw����ux��������c�/��bcj��������R�Xپz��u~/@����<�l�3#�A�����;�.tT8�to��0Ca�����M����k �*�${�yt��k�%�؉�g�Il̜�t�G�،� �֒O0�G���>ʠ�@Kj��xi��
�6$�������D�ݤ`�N���\�,"���]�k�Gla$v�w�~Skj�i���4�O�8_X��\�B�Z,��i���l�����jo��:��3�W>����A�smvQ�O~�K�R�M�.��;)�3C�?���K��H�A���d�;��?���s΃�Ɖr($5�9�i{��0Q�<g|��X�t�"��^�+_)7}C{ߊ�~θ�7�xn���`P�Dy�7K���FGe�	$�Q��K�>&������y�ړ6A�/6LݤQ!iaj����*W`��}Gh�	bьi�?�!6VkL��x+s��%���ڃ��[W����bG��	��D��=H�[���/�/ ��i� ��0�Gt���+c�0UU�~v�[O���f�)*;�2Z��#}�[�U>�T�[�2��Q�Rj�uɫ!�`��h�D:�	4�[/`��A��!W����� 9e <�S�������e��.�]�G��0X�����V�H���4�.���D�C�^s�o���8�͟�����4���q��0+ �X�J&i\d:��i+�#�q�t�J��\:��ܭ;g�[7K�Av�H�~��`Ya$��}�����9�a��O1FM~���w���9��	^���N"s��Op{��3�j
Q�bM���y��]�LV�̉�U�mvI���dp	�c�}��f\4&��:�l��-Z�-��pXz�:�#w�X�=	�����C����H��5:vӳ��v�d�������Y���)\,����$������m�q�.uC S� X�E ��BR�
*�K��#'�$���kKlX�jl��=��i���Q8��<�K�/q%$�·�qտBA�d�p���y��]�}��MH�4���'r�I��§<��-�Y����ZQ$�*ϜK:n��Y.����D���kvB��ih�s�{�o�E)���j�q��
�� �y�	d��0Z�����B*ϭ��o>-6
�!&��m*���Bɔ�`X�v�(3S9_�sx�%���Z?�v��[��hZf�խa����*�1�Ͽ��Ge�$��b�b��Q	ڨ}hQ���ȵp6oJ���6Wr���1|�P�)>��(����t�KYi��٨w�1/��=��قƳp���#T���PK�h��rH=p�Έ�d���l{�f���2������q���3������H�������	���G<��)x�P��|/�VL�Ql�z�ճdG5�ֻ:����t��P��8Z,�}��rҬ�m�4�-���6�1U�e��i&{=����r8��1"�}�8z$�nwL.ؚPqw�ǆ�8%z�Ҋ�@���vFtc�R*��%-<jק^�a���?�-���F�ڧ�\�u]6�/ϖbkD�����Í;Ő�um:҃(�7���J��v��[`�����,�Fe�T)�y�Zi�=�3�p��p�$�Pܽ���4��77�Lx����9[��_�K��(I�&�x�R�|J�N��^$��~.\2�0R(�t'8�SJ��lVj�)t�b��#;�C����ҭix[��ݟ ���#+%.=��@-������'ÅE�E%BV\?�;U������p�Ź	ź�����Ǡ뽏�q�a���d(W1gyqZ_�ʔ�mv�C?���ٯX�#e�P ��ޙ�S�tI0$�4tu����^V78���P7(�8AB\~�I�g�|*HjYK�����$�y�')q��.݈�G!w��(��
�/G�B�����Q���2ÔI�r��!ҿţ���`��d�B��4���s�k8�@
��)vE!|���PEFn��R�ٶ�M�|3)d�Ր@��W w����Џ�ڌKd�*=�vg���ҏ��P��x���(����A����I '��q.���%�p� z)�"� ��σ�r.q.�V���}?�;>�
�i���!
�m�N�~��L;���fJ,�89/��Ęe�y�t;`!���"�jM�׋��1z����O$���2�0�J%cј��$Z��b8�\�W"/�4���ՇDU�ė�"^eP�;�q�����L�z�ꃵ��s�I���� ���`$&)YS��z|�L�x�����@>+$�z���t��@�*u�q��z.�a�m�oj�n��&*Ps=��́�S���LE�~Q\V�J�&P����b�Ҭ(��]Ë}-͡��R.����'B
WQ��!Ɏ����=�d{�&���~7(a�Ƃ���������z�u�RG��.�`r�(�}-h˯l���̤�ة�g��؆���zx�q�kвk���Q�92���ѫ�+̶�#}��~p_��� �b��+gE�Ԇ���o�+���ZA0���{���wr��+����[s���?���U�l);��hFRmvˤ��CJ�KxE;�[J?�
�����7��6]��c� ���T��!́l���O�6����̥�R���,��Ψ�XG�#��|��zM�6wAUz�>/YN��z�\�^�1#)�E��G��&��K��+D��upI#� W.�c]۹d�����N�+ж�秳(Q�b�Y��N��6^�M�\澈D�,���(>�(�HL\�pڸV��;����'��y�(15D��o�\��]x����%ZG%�
5䤥�L�~����H�79�;����� �Hurƥ;�n�� %sQ��ƚ��p^�Q�,[�Ym�ċ��sʬ&L!;�����oS.�zo2|	ҏfZ�s3�)�1n���)�Yc/��h��+�jE ����-L/pXlxVHYEB    fa00    11c0�iL=��G�mэ*�x1���F
�x�
�c�����*�E)l�(܎�z(����Kf"b�g��$qy�<Ҁ�K�&�k���\���J3�y]Ǆ�9�����-�Sm�ŗ>M-�q�C��(�}�	�� Z�����F�����W����u�6��EH)�a���}�p��	8j5Ț�j�?3v��p(�>:�E�Q�jZ�*A��/\����PZ�Ϟ�^��{г��َ�!����W'�̰(v m8u:Y�� Qz�+��ٙf�*��-/t��xz������M��6l�W6��!\�A탗F����Y����п�JiN-�<��$��z�[T�aut��|M�-�*]q>�"�;�)P��3R��A\��$�m�򬫥�m4E�"���?7&�%�8��)�a����l����&U�P���5�U�G�%���
�W���+����%K�ìd�Sf� B ����-h���1y�� ��2Gt#Nf��Z
�����6����a�!?7_�5yʗ�݌�m���R�������hI'��Mx*J����]{]f�'q�DW��_,�Gݧ8�W�i�@#���`&�Bz����j�/�49���b}�S��$W��IN���az��� _���?�h��73�� �/v}��10yXm�"���oHS>�vf,�G��X�w� 8�ov��03cf�{r&Rb-s��Ƭ$��Q��B3OmSVb�B:t�8 �i{5@�|/hʜ�r[:&^b֑����Peɘػ��k6��9����_��v����J��JC�&��D���A��ϻ���jJ]A��7k`�_sy$�6�������L/���H���ŗ�I�ҽ1�.��!��K���L}|Ʀ��q�m�j�^t��!�d��7>#�"��i�o!��sls���� ���Ӽ���<�׺Ns�o��8Ɲt�Ol��tgm��n5� �,Ks����m�%&��[�1��N>��S�˅��16>�GS&��RX��t-(��%�=�K�W�� ��'�M���ݽo�c�41�hc<+�[���A���������1���X����;�R�Q��n��t7����>Pb(v4���F P7�}��q*�җ��8Z���?�Y�Y6t�S#zCQ��p����w��.f�T�@]���4C0>(��-v%:���Z�#�\�eB3R��"�*Y;1���8���/�REk �̔�'o�>��4wp ���L�)�M=�� ��y��S�3��X���h�0$�cg�c�,���6Pм���
�|G�v�@Qyai��n�v�[�x�VK�kQ1S�KK��^�{h�b����s{�x/E]�;���p��I����0�������{��!w�3]P�+����-�WvŝF�`�}�5&���J_V*|��o��IJ���� dܛJ��S@SJ>�	�0��q����Q�6��7���|S�<2}c�۪43�M��<sD�q<k
��!dF��g�_�ءG%C���?ii��x�c���lX�>�w����2�M��	J2�^,vJv҂"�j��v^S�](K�Q���qu~9���L/�P���Kd=��fԫ<%�i8�3�ݒj0���-6�%}�[�0��΄�����<:���ڠD�z���e�����N�Ld��NML_qBJ}#;�#f�-%d�H}h�#
ЖQ9jv�T��T�tƲ�4���%�5�����X�Q�Kp��sq��O�sg�����	(�����g,�Ϭ�S�
�����G\W'Oaf[����)q�ʤ��ly�L�|�{�Ň��k�}�w]�w~��Q�_�dK4��'S0���!��z�b�|K�X5�y�b������Q��YL�so^�%���$�8�մ�XyΝ�:��h��r]̂J��U��띨��c�Z�(厾����"�d����D���ir��Y��k+���ur���O�)O:)M$�J�� �֋Z.�c4���A6n��ڛT��^u_}��F"��/��B�K�o�X����l��0w{Ӓ��@��8Il3�ԩd-����.A�I\LA�A��>���_�)5ܙ,����"���`���H���Z�������4|;oG)���!�`|rdCs���K'M����Ö����G!]Ě�+�F�޽��_�-WkRI�33�/S��S������Z�����0����罜�PW9� ������s#$9{��w��'_��C)�)��(�W�Z�<�Z���,Ŀ�g��h-sʈM�\|[-{�ŝƼ4�.�g��w�cD�\�I��Z�|��x��cC�du��s��/n )�'�5o��`t��n{	Y�����\��T��1|��LA�n��`[��d�����di�z��{���0%M� Y�1�s�����5՞$�o�22���1kY*������N460�����$��Gݥ3ykV������6 6�"�bR%O��P�j���bўYU�n �����?�\ȷDQ��=|"�Ƣ� m9�*]��.u{3$��a�kʯ$��O�O������th���8���%�r��`,��k�-�����Zn)Y����!����~��\��>����&y�nޑO¤��d��y���Z��BNG�#�@��Uѷ������2j�� |�"��_�j$K,y�^��E���9��؜�%���#����6EI�y���\�?�g[9X�bP��g0��Y���y���8U�f;�2�s��U�f�Rh?�L�/4�a9g���N�T�L�"ʾ�H�'���Eg�����%NIR�	1k�tI�(����=l�m�1@� s�9�������m!��.��H��b�U��)bg��M+�a�%�-x�	��)�{�WL��������zǣ���C��i��L?GQ7$��O �tYQ:4Q%�L�P���M(�\j@��JB�uԇl��l�$��Kq�CSخM�i�^��fy˖��F���u6�w>�4^�؁�mt�5�a{ǹC/�D0�ѐh��o�YG��Q��D��[�~5ZGq'8�t�7�E�O�+B]i.�߫��BCi��=ԻL��|�T�E�~j�@����-��lW�ʛ;��x�BN���ru�����l�?�[���v[�ގ�("O��)8�W�Az�S�v�ON�<��H&V��>�U[���"�`�V1g�����/ �e^��}VBNߨ��D������j1�(�?�D��^�u~��;�k��Kxl��� ����J�[�f5ה�ʁ�\x�ZN���Q�����)%�!���u�+�sF��
\u���2���"�����G��	eݟ�e��Bs$�
�9��Kx#�H�۬K8�b�v�{�n��UR�܀փ�����������=8(� �`��h�7Uv�s��N�����sI2Έʗu��Uy�WW��I�^�pse���'��cY���V� �X�y�C�{g���)=u�A�~ߖ���V����=��8,�j���9 �Z��ӭj���@��de���Č�C���C"��9�>�&k�Ж��'�G2��kRhR��w��O��6pFΣ�LJ�y����"ӝ��%�۠�o���w�^6�+��2�`[@�,|$�q�j{�5S�g!745Q)	�Δ�
T���|T:�cx9]1��T����Y��>*.��ɦ�.��A��67`e"�o
K3v矓���k���y+��I���V��dV딿��?pgjXL=��R2�[G�����ïN8H��P1`�]�Û�Ǎˤ�ec'�ԹM����A���W'>��Spj9��L��>.	���1O%6�љ\c�E����hi�y�	��zlM6.�`'�/�]���w}�"	4�M-�ݐ��=�
�r&WA�x��,���1LX��|���/�A�n�-����K Q��m�Vg���2OSܱ]��2�I>JD�;��N;X�˪
����T�|n@)��ޠ�ʡ�j�]��� ��?�;w&�<~�~����b^�g_��/��YL^�Z=I�����V*���p�~�5�~��o�n�-�pO��/��H%�L:�h,+>{�c%��@�ʷl58v��%�Y���෯1չ)��E;�Y��ɝwU��\�ĳr�[;r�ʭdn!Q����bJ����%F�w.�LC{Òv�*?��u[ϣQ��|
�^:n6��z�k#�aft��ܘu�: BFz�!��$��1�+���ud#�|ĵu�������G���9��3���nZ��+������E�T-��!r����as�ɪ<@؅�}��cS�2���!-+��*�csP k� (>q��8jX��5���6_�ͣz�++I◻zhv����~i���1P��~hk��Z\^E�d��kX�ލ��Q�G��WE�PB�RZw�	���l�[�XlxVHYEB    fa00    2cf08#d>/~��&�7j;=���6Z�{��T���_�w!���7Ct���j΄�����E�"=u6άm�*���ȖMxI�GN4Ll���Uz��� �O�=S�A���Ɗws��v�u�uh�h(���(�#R> ��wtnv+cd�9�3Zn#V���Q�Lz�n��hz ��C�՝ y�7%v�vS��"R��C�B�ֵ�0
IP/:v �s�.Ggհ�t��������c���a�IZ�'o����k�"�&�A�q0�^�
A3h�hx'(9E��L�v�!^�L��j`p����<�q�l��!@�F����P���b"^��3�����z�*�z��/���֓��y���?D���]����=�-?D��A֥�FU���M?Mؤ ��2*�A�Ԯ���(�Kn6Q�|cD/�+��ӕu�h(=N剥mR�&?�1o���:Q4�E����Apd�ɛ������H��od�m\q��B���!�=J0�$��n��- '�_�(��"B���N	&�|2Y���
[Ĭ)&5�/�34ϥn����&��[(��B�/� ��J�ޱ���q+�9���n8�t�p�����u����3{��c �pf^~�"K�W1�d��<ފS6+��>����в���FN�������A��|_L|�,X���[ 2sO�=ˊ.��$->����g2L�R	]�u�t���m@�Ê����1[�}`�>n�{Li���t�!YM��*X�(=�q���"Rҕy�"���V�H��B� ����Ĝ�֫tc��w!@4q�O�WQ�ޔ���˻�C��ML9S�o���p7ج����dH�D�w�Op�e����\Z�l�e��Ί��
_]/��I�a~@�A7�/�]yX�L��j�#�.^Y$d�hğ��hl��ݰھ+
�Qʓ1繉/�]��S��<�"�\�l�ϋ�Zk�4J�����/�A#/kVhF�/��o����^u���.�R� �d��P&!���Á�t�k\~�`#C g�YkIBb��-��7p�BN{����hz��ڙ��r���P9	Ҹ4�C,VJv(F��O�WG��na%��LƽĜ�!N�>�Lr��)J�f�=����b|R�������l~Sq�N��e���C3�"U}���秾V��E���W,H�����D�K����B>�v�-�Q���>n�(	X���`�F�t����pi�E�${˻��_�e	O�;��AɄÿ�M���B���'�"��HY*���S5C�[��[��E��|9dr�"�r�vlh��1��a�b�&h�bi{�<�TT�A�|)7C���#�($ G�D��7�v���_�Z�rW�͘~��.xa <$�*1d
>$��ԫ�ے����M��O����_��>�i�g�����N�rv����Ş�/�����fz6��Tp�Y����p���>���B��ĉq�a�|���!��M��
i`��m���z����'l�ŜU ;�}c	����t�q�L
���&0a�Կ����Zm�6�~��i�(t
g=R�辕DM��$�N|�-��l�y$��A*p��f�ߵ�̾Îr�G��JЪDV�I���6�u8��`e�M������w� .�+UI��y�*�9�]�IkQ;a�b����{��8:@��Y��K^!a�GԙU�i�(�&udW����CKW���u0����n=�>�	����s�ozckX^�{�φ�����[�u�4�����"02�B�x��3��bET�x�ev ����o��ud��EM$\��H���ԃ"5�|{�L�S�狜)A����\~��`i^��=i ��B�>|����7x&"��t�2��F�O)��pD�k�s�[�vI,�b�U�3i)�U��"C��1��
�֖qm���љ������l�UX�������[�����H�i��e:��WHtB��d4�{����ҩ��u?��	+s�ҍH=��ߎ�NKF�4x��u�^QWe�R#��W��EIrpG�N�a�As���`�8JZ%�-��?�v"Hp���ñ���C��Z���֕Y>��zY�s�����`�>F�[�b]�i�1��M\�R�}�8����]��Ah�ϙ��`9�'�`�%YX�mB7����c��+��8h 5<8u���T_�����Y���6�����nS�,�Xo>k��Z���r�ı��d���h���.=�P8���o��vy�@��4(�Gp5��^�~�]�� ��!r/4Ʊ�*���qÿ� ���Zc�A���6�c�n��������BY,�|e$z\�3�$QI�*��Fg:�JX=w��l���Λ0�����P��ٌn����3��k�U��R��3Lg?�b�Ue����/���$|Cd�!خ
E'"9z�j�i�r����`FXXbc�?�_HOl�l�wYcD:�/N��	�p�xt��A�l;��gWc��D/�-��s�[ѝ{-w�HK��-ʳ�u�ل�v>}�|1��F�Z�%#mHh)�f��3�������������E@H2$��󐹥t0��5��N0t;��^��ơ��V��(j5��!>,�"m��V�j��y��*���A�C�V�DG��E����HA+��Mj��qXY��v��f׌�rE\Wj���!%�������`�}�f7p�Ⱥ�?���w#�R;|��T��J�iwv���Hj���H��p*�eX����hqJv_�$.�h��.-�T.y�]pm��.�1��߬]U!��ɾ��Ů�S�[����������l,��Lm��7.���.D1�q&�P�ʈXn �� ҃�J�ڨ��p�ฬݘ�����j��3���Z>&\���2�x6w��t�l�:'ޝ!nc_'_� �^�HA����5ׂK�ևv�-+�����}��	��OB�qbG����|������R:T5�S�l���\F����S>y\��m+���d=�����7�}�y�ì�@!���}	mxW��X�@5��~�G�}_��%=��rM����} V(�y���R�����lȽ��f�LX��|/�Q�-s_�"F𽿛l�u���K�ŕ�¡��A��
�;@��IT:�z�H�]-P�>WLY�k�1>��eA$�7�ߓ��/���O�sH�q��.��m܄ު5�{z�>� ���� qr�Ǿ��I:�\�|}}TC��S�s�?��DRo�{%&��|v9��۵����F*ׂ�U�a�W!<[dNU�����=ki4�[��,�3�
g�O�	x��&�)oE�T��?\����̲�X�΃E�zө3%yE5��Z���9��1��e���-�1UgƧ�X`�L�}++��R�m9���-Z;-����z �"�5AM�0�F>qv����ݼ�����-�-XS�%���T_N�B���F�7*
�X�/9� �օ�O����1�����--=�%B����܊���v����ex���%m"� ���f��#���Z�t�PBL�r�����m� <AQ�=���鸦3E1OruTa�$�B�	�'��=<T~�t�����}r�H�Z�f3_��d$���N�9'�d*`
��O���'���h����_۵�#��K^v�B����O�v��f��̣;�h�m�4Q��-E��{��ȑc�W��LU�� �� e���#�>����6��S��[��$���O#L�L�8�6����� ���W�O��6j/�"���(��Q���G�8���4?"<�vh�����p��;Ic�a�mdA��g��&��ԑ4!n��0��b�<�9p��c9��U/��):�Q&kxj���H�#%�fɌ�Z�� ��Jm^��u@]$�(%+���o.}���K�M�kWXsT�%���]�qv���m�c0��!�	H ��N�AMip�۳+�N��pq���nc��S����͜��Ƥ�}�3�9�_$@t8n�h�Ҍ���z�yRAe�����͂Mq�Q�?HԊ���O$�
|�W0	�І��ʅ�F/Q�`լ4��^�r���$�6��<˽%oGJ�o� �w܏#������e�Q��xK�c��.Un*�?Y��kkm�d��m�{'e c��PJ=�����7:˻:mLՉ����#I��X�ڊ:��?�,�PL<�yZ+r���<�ۺ�5r{�RR���Z$��4��*��9R.��=�K��P�mXL>&M8PYģ��c���ɪQ�Ak��@@#+�E��@�hue�'@YwJ2� ɱ���8^i���ں���h�cj~ٷs�����X0�����X��>��6�T�o��aT�a�Pl�s�^� P�`��+R�{���赗Y�C.�k��$��$m�R�#'o" ��F�%T$u:�����a��k�������Iu\���4�y8V�@ЙHٽ��`Z~t�ġ Z.�:��J�`��d���T�[��s��+�����������љU��@Vנ�%�1&E�~Q>�������_�������5��xhP3���咢X���z��ң�T��N��������������rU���ӡq�X�tĂ!r"\�U����=�>Y�^�.�2�<������)��"U����c	ҽL�c�W,�l�O/K��t�^X�͓����K4]M�bl���r����/��І)��,J8�S����[Ny���_�T^%�>���"���C���J�W������R�d�}��F�1 �!���N��
�z�+�Q�i��i���){.�����R?l,Aq�%�}w+���#��vD�LX�}�{Se�l'����kE1����8�=E�E(�G�E��e)釕�������z���{��ג�$�����"%�����Ӵ}̣���#G����y]�Lq��S6X�׍#�~�F��κ�� e����&�y?na�JFn��-�I�)�y��ӹ�Լ�)�E:���??r*�pg1�r
H��E�C���I-%]Vl4$�_3->�[Ԅ���b����>���8b���a��Ni8=�ѸJ%v���6�D��� �'�r�����/�Y�ѵ/A��m6�1l�#��|��bg|'�B�mV�E�/�Q_�Q)"�g^�Et4��S����5]�q�� a��G�������疯
o�<��X(�Y���ʁ	�k�C`sd(�A���	^]u��)2'���;A�X�k�`V~K?>���hHZ�2�X��h��t�W�0n���H@@�3�h��r_���k|��h�Fh=K)��Z��u��"��(��+M'{��8J��i̟:�]͋��C�l����#nB��eg��=S���/���Nƺ��U&��}Ȁ�f���G�`�I��ֈ����`ۦF�z���H�7��R�c��[qsJ�X�����`����N^epL.�I	dN�rr�Q>Mvj�u�I��0������w�Eu�2�p��F��l՚�rx�2�8{b�"F�+}�u>�)5�@�K�"��{�j�S)�@�/����Q�F� :�����n�?�/|k����`�J1��0�][/$�$T������n(�����G��ChJ�X�'W��2�<L[�u��P]��<}��;%�&N�k�n��9Q���م��������m���r�$Jେ�rk`NQ��(�gZ�j�� 0�����Ȭ�i��O�v���sA�4
|�E0�`cS�i�1�T�N ����Z�*����q�����w��E��|�N����ҋbDl��T��w>�&�r�J�\ʄ��"Id�* �MC��\���P�"(v.Y[���Co��As6n1� n��~���h2󽇤V����b��BQ0k�aZ������*�f�z>��/���H��ܽ�^<1җ�|���?o��~ Vf��I��k�g��m��M�g����E��R`-󹩱3M2鶢�
�R]H|�-�CX�ӿ�H��hh�NC����xGu��gT���[y�U*��V�O�;��VL�ۚ��2a��e�$��e�6�?��Ge��=bp���{�_<�<��}��"@46y���ވ�+Tf�s�tD�^��[������Bv:�z��] E��}�UVZ�n$�Pb��{}WOv�G��g_� & ^�tj�2O,�%}�w�Bs����af�1m�^P~3�r��P��V!��#���ٕ����͒���[GD����`���,�8K�â��(����:��7T� �jJ���҉�v��;*3L��Q�D�uu0�ƺ����1�(�#��є�mIRs�e�VKӲ�D��-�u]'I�ӿ&n��%�h�~A��4�d��@��UcȬv��K�Io�E��ôy�{ࣈ��s����#�l����(H�5D�L�y�����*�(��7�oy^K�b|�����~t>lX�����:RØ�W7>�,Ni�,�y�,~�fh���:	��a.$��ф�E�7x�g�B���{#@s�cy�َў怰�^�cJ!:R$����U���L���#SO4�,qA�=���W�o�W����&�xh_��������͊Uy�I��G%��D���!Ya�Uo^	E��R$!��� �p�8��N��rb_WI2L�՜�a��;��^�"k�/�|WA-��u�"�^���S�y�OC/ss�w+��'u�=�2�̘o���to�X5%��FT�v�Ј���HT ci&�W��&JGq�WMe�-;rC<�T� v_��y&���}��(5��)�����o�}f��^�B`�O��4x ���O��%�~3��@[�A`Ƌ�1���sj�_ͤ@r	�н�^qq{[��0�nc���ͿL�����K2����fiyXS��J�?��w!Í��~� k$��ǟ�F���MY��8��̖�)�����D"�<'�U���]��W�/�[V��\]����� �AD�xt�b��3��+,�J�R)e�O��|�|����g,����%��t�p�Ȭ�'�׀u��Y �$��.�7��,'U�2���̸�J([� ����-��P{d��w]P��qę�C�f��;:���G��&��?��{95k��s�sSG�nK�ں���B&��L\�D��pꨭ,�ʎ�W���Q=�y��'�
�IX���gFCj�ROy\����ft�����o���zw�PXҌD?il|��x���Gs����s�!��'<��a��=˹2������Ҁl�eV`����A_���'�rm� ����&�L�O>\�Ŭ���!��>cq9�կ�2���%t<7�U�J)*pV���g���0e����؅jqM��x��K�^��'K�)W�fAA*v �[!�o�� �;c�O��N�x1�d]@3����XKUb�C*���^D�u��:�R�u�!,���\(�@bqNs�m\�����=b�jtO1����ڨ^�f�w[�H���@�a���t`���l��W��e�ʋ��R�[>▢���5��������C��9UA)<�`=Rs�.Hi�s�|�P	�R`�R<꫉N��K^$�ey���*M�f\8�ߞ��i��^�9�y��N���m�z�^�l�y?�V3I~M����5yh���Wc �m��B,�djU��QL�;���;�V�I?�7 ~-�! vgm+�.�ho4�츌��L� ���=�;��
��9u	̶�Z�w`�;���M&ǚ���>;��d�
xd�q�҅BҞ�۽��aґ� f�)����B��>G<�����+�,�
1�;�*s^���WT�0�`�5-9Ξ �q�����[[�Ƈt�[��z�ZG�a����h����p�̯�@�`�Ӵ�8��i6��g�_��Qە�017�9r&F�=��u-#�-�G`1�c�=�%E���;��$K�vE4�(s�T���Ӄ����M�Gio��p� I��{��M���U��\���-HT�y�lP�Ѝ}�sd�́9�*zrp��\��^F�k{�S ���o#��$�1�����7�[?%,	�beI�uV+�������2����hl-����r�^xtpt��I+~�Np�.�P`T;�����?��Sݵ�d�s9mٟ0=�?#MA��v�t0(�bSz�����Ҙq�~�s6�J��_�o��f(�uow�\�$.�� �j����ŏ˶ ;��#��P��>�2
�6m~K�y�#��kЅ�տ��[w�!�w��c2�?��W��$\Ӏ��T��e�_:9�{���\r˦az���7x��_C�)3�z
����WNڗ�u�/*�v����H� �KQy�`�A	�X´Z�F�g�{�:���|�s�`D�^A}yaL�-Sf�c��s��h��L2��@e.���箺�)$u��e��Pͺ.xO�@|$+���P���?��E�S�^�]��#urL5�±lo}rҴ��S±��ĉ���|�e_"�=���̋X�bt2&!k����b��qV�����?�C���k��<��7{�}�iW�uV��4����e>%= `�6: �O����Km��k��Q}�����O�9U��kh_^L��R��*$4�a��o��!�;qOQ:���.
���{��:
A�0�5*�l���
ƶ��;N5R�x�8���� ̏��7�)��a�35;K�rR2B*iF>��v���el��ṟWmq���m+�Y/C�M��]���|�R�k6�ŧ��{�`�i�]�@��%,S���*>l��a����Bx��vĲ�3�/)<S�s��c�ңk�t3\��h�oD���<������';�V�4�]QA����ǩ�IQ����gfkˋ�.��%��ׁk�����T�K�I�wuԧ�I J�'w'��`=��?y�O� ��--�s���8%�|z���&���-�\����Q�S" ���r
y}�\W`��ݕxK� ��(��th�g�3 J�5�!*��-���̐�]B�Z����,y?	%���86�C;X,��$�A�?��V��#e}��c�xIc}u�Y�q�6�>غiصm��I��/���O�U0�=H�����糨0B7ׅ���8���pj�'�*��Wl9��e��{�aE��z�5����q����Ћ���NG{��@T��T�j����g�q�ﱳ76�)tk�¾�J�rۓvzO��?s*%�9ǿ��l��3/A�F�h���b���"l!@����>�5�����/�)\��Tľ�Y'��
���Ҁ�>d��}n��q����(~b#~�@fS��O��;�ڮ�4:�ħ����z����Z@+�ا`��;l{(�ӓ��^{�j�T$�������4�	���O��V���+�ؒ9!�M���=o����{�y�����hJ�ќ�i�(]:��8��e<^�_��)�`�Y7�QX�Q�OC����Br�u�I����#����� �
N=�e���%-���8���-�FA�n�9�}�=��M7+ry_��b�.b���&�)��ܩd���	wH?��z�����B����f��o8c��X���:��X��`��gxN-r�����qe�G��t���iA�_,t7�vRH��R'�^❋�$7cˉ�Ĵ��Ӥ<���1�S9,خ��D,L�<<H1\9�R���d\�0��q�x�����e|B �2q ���2yf('a?������Z�>��I2=�j��v�8���з�V/.�W�+�`���iJ�2m�ċ����,�m�۞ܫ������IW��Q��(ǚ�}
����#V\�IN �z��<���_�4V	���� �#ْ�!Ƞ�S�i�o��GT��h0H�t�ڐS����O8�A���0���B~ml�lF1H�>]��`_D9�E��r��P�Q����h�}����x\��A�Zo�_E'�K��PG��yn���+&T3bh��/�]��v�b��P ^��JP�݂�#��f.�29��o��tC_���8�2�E������>OѦuߎ����U���v������-f� �Y��/���M7�,H\�Ѽ��kNe`'�ȱ���Y�}�~�iLlO�(�h���V��C�v�&'��7��9B����d%�7b˹Pw�¦��0o��Gd�܌�u����PŦ������X�7?B�V_#�sS5>��ͧʻK�ʏcg�:�yRDRHq�:�g�����@��i55PM]U��B�� `��PIo��_s�($΅j�HB�1���2|�Gy�8�1�(��\�r�i%�튜�ß�Pʆ���ym>5�gq�~�k�^�!�,��a��)\e���g@�G5?�$
Y����vlL��늫kK�-V�p�׾ �H�9ըǞ�<j�A0��g�Sv`���Q}���3�	�r�������*�q�t�n��㗕�a�cɍ�l�.���7g0�jt���6H��j,���PP�pa����j���	�g���Oz���d�͊i�*��M^R>��{V/QF�mHɗ3W�l>�t�x$)Yr����w�����ܦ�͐��;1�x ��G�IgB��rJ+�Ș��}���J���;F^"�]Sv��|�1���[��@����?��H���l���B�*C��&�¾
�m�O��1Fs"n�9�v���J�-���kj��[Hn*&ʾ:��"A	�N?����4�ｃ���fGmU#kI��l��|A�^}��`#���y`�X��Dj�S=�+� U��ꯍ&�7��{�Ojb4�a�'�M9j�!vS	񫷺���K��u'�l^��� ��g��R�'�C!�AizP���/V�5\z��_/$H
*pu͟�i�8,j�����g��N��������Ld�Q����m���ˏEu�Y[�r���lU��G��`�M��O`x)�I���Yp/�0(��G:Ap?�c�o]5-�K~�y.�v(g��mB	ŝ���j	x���l@�Ʉ.��ÕZ�N"�UA��W��W Z��𐟥�P����� ��<`�@OÙ��9�4�����KG�F�P��E�3�*������ҽ���*v�Y��? ����کd���k���.! W�A�]���v�������;����[�]�z1o2��O�(ͤ��Fy����BN��@�[�y��7y4��M���T��}�{�D��Pt�����f�^%{,3Gm��K�ڊ��^����W2��*�jC�e��u��[��������q��;�(��w���s�紨�MW�˕�0-f(�K�:�/VH\�'�R��l;l	ʈ>.�����$���@|9�F*���g�Es���ͭXlxVHYEB    fa00    1f60嫳l�&�
���޵�o@k�� x'�4��2�����-������+6�Z��ɑ���:��q��+4,z��P�ˎ1;�$��̊��U���+=	�l�����l�ow�Q{}��:�y�~���E֜�=*��KC�{��,�����*e�3�~.���?�0�� �Ȣ���/��qB�B{���89[�bͺǨ���[�8cs`n�Ϊ���-��%���.�~em�(fR\��*��������K��e����{��`'uc�z� ������h�j84ͥ,���
�f�/�`XF��˒<3�9E<v�'f!��*�k=Ǐ���7��F����4p�P9����dڜY��wS8�\�\����.�.G~��L�J�Y�5�x_������t�~as3�p�����������,�8RMll�v���������!Mf[����������,�+����'��[-�k�I��YK;������t��3ؤ��߷B��{��'���I�|��g��P�q���z�j��Mu^�Oj&^��̶�u8޼��qՁ�u�i�I���X���)�9�?Cj(�͡EK������{�a �����f�,
��n]���#*��<*}��q�: ����~�L�m�����GL�Y~jn�`j���fa'f�d�_zKf�'G�I����yP�{~s�YIԵ/�������_3vQ:�g�B�7�'<zY$�/p�~�0��K��l�R�a� �J�r�����`U�0����~b����l��h��M��N���t�ѯA�>ł�\��f12�^����,LY�ݽ�H/��2��$9��^�(�1�Zܒ�FW;�%��I��pO��E\�O\�ͼ��_�.��r2�cF�z�5�/�G��H���w�1&WA�c8��^	�*��_ �a����C�����_�����yO}�]���I�Tv�y)	S�޶Lo?��:��r9L�J�|=�?�}�'�-O�9���T�Q5�K3:���W�8�nX��\�Y=*�u)ԐҘ�� Q�-cχ{�`xzV������GMT���;���\"�������2���?�cfU���;1��ç���I/8��Vǟ��rX�MӍ�ǘ�XM���TA�Hn��ﴴ��=�R	�c�g~_��LV�uB��7��&����W�`�y�9�:s�n@*:M��� �au�٧�[4�}IAE��?Z,u�V��M|�O�yex��ħ_N�lxX�~8{��ηd���<������� �
e6).��Z���uo��qQ�%�<~�����h5m�,�Ń�N�<�4�t� =c��59��`��
*������ɏs:������u����̜7F>,�����I-i)�t�u�z￪-F�����& �q�}�'�շ���A|`�	T�h���`A��=��O��k���zP(��w���x���J̽]u�܇��g���*��s��\�&�:h�>��j�]~�"!���3�8���iw�Q��!��h�mAE|[���(H�XtI�y��[�6a{��]���f�C���?���:�B�c�D�(E���m �'����[�]�MԐ���@x��%薋�ⶒ��\�Ms��g)]Q���'�)�� /T:7\��x�m ���'4c"DAi�,�$P����g/ɖV��ȧOW����&
T�B�zc�U:�>:�����y5�$s���U%Hs���l��fY�|�/&�X����*.�b;ml?>�{����bl�g���-�3Y���[i��5$S��2i*��WM�I��e{
(�A��:���\���F2��I����|@�j���OÃX[JJ�[�IX�} �5�����/�/V����ފ֕�؅���I��nڹ.fVw�xA3�Gv�v�V������J�+'�q�VJ�ZU�â1nl���0ڰ�^����Y��Ά�S��iW �V��N�j��x� t�����-]!6pר>���R�Q��C�diL���"��������L��+9�B,� �"��.\L���IV�>�9��>kD�ܷ���edS��Ƒ��J:���2�Ѕv�v.{�ײ'l����kZ}������-�9�`ʕ��ȃ���7!�@�V�m�u-)ʢ�N_8[��bO�����>R+^Gv�*�Ȼk0>�sFj�̿e���п(�n壝����<�L4��첚���'�Õ���-�������idex�@��Cm�K���cm�y���dR�X�h��k�|�j�	|� @�&Н�m��Se�@Ӽl�̹���q(��d�JV�5�;�xhV�3�����l�l�RC��z�=�**+� ���H�Bd��n2�e�׍�1��$1�,���:}�L(�K�}g�`9�;t����5���L|c�܌�.X-�h����5V,��6��%D��� ��[�^8�MA�E%��>d|B5}��k���p?Px�§	h��8��,�S�����EH���Z!"V���c���I	n��7gM�P�\ *�X �1�o.+����d��6QG��)7�i����W����<����U�Fr>�B!!8e����G[�U$�Z4�T�Ρ@�����W���q�*��SY�\��{F�s���5�Qb؟ ���E��sl�$s�N��~�$��C�1d�ƀ��oK�qYF��[��[�I��-�VQ�V������!:�~^���̉�S��ѐpRݽ\���x�ZYcO=a�N�Qvu���f�w%�x:��QL��^�]�
�� ���l�	E�1>d$,�:��/ȶC��4�i����2��'g,�h�W�t�H�����
�S1�mUg��=i��V,�?j�o6Ɉ�."5�u	�Ɓ&C��K�e��rD	gX%����n�`&獄�g�gf�2s� ����NŷAY$ą>Ia7c����O�EP��s,���T���T�|v7<�tR�7��crd�����'R�".���0��#W��4�)���)�B�����q�
�,�]O���ّZ����B��3���K�i���	Cs�Б0"3p&����}��FA	���YA�G�A����Ӡ�IM�IaMP*��%�z��u;G�{��N)r�A*AlF���+8��e����:r $h��A�s��2=��d�
�d���_�K��� <Uk�.]NH��Y�n���e֕��������"���.�%�BBp��uA��`J�u�ᗙ�aLNQ*�������R���\H7;�a�A��]R�w	`��	���B�ɺ$M�گ�/�@qc5��@��R����W)��l�^8
]�땗��J�����G$����t��[˯l��^�t��i�E��Y��k��וwj��EO���K�$[��Z�|��p%����e�pE�>W(`�۔�)�k�Y��R�<���8q��;zr�5"��f\���a����s)��5�V���D]��w)p�'9�qo~x=��z1����uH�WU�)���p��j��ٶ $(I9%f+��;o�ij����$d6���r���bI���WF+�Lˊ>(E�#S1r#�#z��]Bk*�w�|gr����0��6�� -I��/���d}�R�(w���ǘ�P��w�v��d�mv�@ T�[���Kh	�Fa���O�dć��]�J��>a(�~'G�����"n�w��6-�JTe��>Ppqy���k���V&�*� ŷ���b�v!i������mHF�2�D�F�=�pQ��)�^F;�6�F����<���ZNOj#W�	��=�BZ��}Ҕ����˗����I.>��V>��Ϭ!�%��W�N����F/Q#��2=�³ �����E��Ugg��6˓x���<]�H$�<o���ݬ�zO.2s���'sM? p>x8�l7Ø@�{�d�I�j�Z7�I�E�m�6�Y4�@.��I���Z⋃T&��V2�2\:����i9��S�Q�f3�XTA��j��]��ʐ��y����/�h�⢫�6қ<黇��<������D�ء��0�.��
���
ߤ�����7������b�}�C�Ǘۛ&y�NE��>�IS̸�H�ә���ظ����?8q�eH�$DC6@1>�;�z�6�vߺ��Xԝ���D��c44~t���V�r~�nAn7� ��S)�a9}�BL�F��h,GGV58����Φ�h��;P��w!J�q�4W�����U϶*����{^ N7�IkW���9_��1���nu8��>:o);7�;�d\'��m�Ϟ�(�]me�����]���E��hH�r_g\��¿`4CfW/5�y!��y�(v�G��9Ɣ[�}]���Z�{d��2��<&Rp���gcS���<?q�Mҁ?�M�e��l���01:�L\c떗������5.-�>�;�)I�M/P�/���3�:�x����	4�幡�r~
���+�
R�n�Ch�[ۨ&2�ޤ�i�	��o���Aϓ�{��O�9W_�����	٦�~%E@)�I��S�j�
I�&:�8��>A�����}E��۵}5k�=��4��W��l���X��|E5�Q�ݦ����d�%r�9��5I�_��qH�����l&1�3�/��xZkϏ�v��`��_bM̀3��z-S��X��@q|��.�h�����ZTF���V�Djp"$�Ƒ/4m�^m��.��8]����mh?�ߏ�f'U��arH��]����Ct����ΕK�̟�ei��3�)�[sx�i��2�mt�
��+@ǭ�H�u�Gm�W�H���z7�xrr���xM�����yY@�*���F�w���
�an�u���ʳ0���)1��
c>���#�^9 �9˗�Y�ƛh��x��h"}�مYH�� ������ꧡ_=�����=����a�Q�91���`DQ����(=Fʚ<�o����c�L�.{k���:˅����\��J�İedZ��Gu6�޲R�Gꄥ[f�3��|	�~W)0���H��Zar\C�hUZ�&�Ló�+�߸5���8-�"�-E�NQ�a�7�\!L4��ʜ��$K��w-��C����:.5��pN��T^D{��ĩc�T3����s;��HʊƖ�Uҡޟ���������+H(ۅ:Mm� C��3��D&�>�zl���v.l8�gt[9731V:Z-d��<���@�!9�(N�[�$6��D����˧�`��j��Q�XHZQ�C�,v���7̛���Ǫ1ٕ<�,�j�8܇��o�����&1N�q}�gSq��� ��)�cK�&]Y�q��e��ݷ����TR�>Ք�uX3;R�޲��z:=�gV�!Ŵ�}�WdzI��[i�߾��#_�Hz��ܐ�?�@���?
�<�?J���X�Eh�V�������q����F<э9�j�Ql�gB�ӽ�S�Z�ざҷ�}�	�܃(�M>��8�Bw�
��Qw6X�\F)<��a����2O�����M�ᒺ�+�y������k���9��\Spg��ʉ.Q�#�>HI�n����s�[?���u��*�����QZ:��s�D��7��	��j~��詰��r�$��e����|�e�S��d�c �� !ä~��ý��+���ét��75/y~�M����9He" c�E�賨fE�b�
@]���8>�$/�ܳ�T�2�pq�V}�񵒲t�H,�c����
)0�iG�����][V��١(P0��������k8�P��C X��lTֽ[��������k��*NӪ�%KE��=��c1�v���|g�M�>�ס(��`�jeF�rA�1�Ba���(y�/��_���#��6ת�V�,��]�ox��n:�W�-�6E��9�z��&�s��f:�Fw��%��*ddo���^����0O�@{m4Zs�O�O�ǰ��4<�ɶ�i�5�ai���{�{V��G�ʈ�z���kfы��0�O���Ē!�~ӄ�R�l�����猩g}}�>�}\T��l@��Q��L�~��W�Y+��� �̇����$i'���Ӄ�u���h݃�
.2��2�
���4i��(�[ɖ����Sj��5��^�2=�������|��c�>�^�Maq4�]��:L��H�ȉFx�KNՅɪ5�+�pG6�l:�0`��X��ȫ���F�=�~�0��m�P�d_-�E\$4��ߨo)���)��H�MC/
����k����f�B�:(+8Q��i��&�.��e�ܑ�!�O���`��n�������D��Q�?��!��ֿ���kނ߁zG��wt����ym�v�LZ��F�r�]KڬXFi~)#���x�6R��#W8�!3�p�	���{�Eȗ����~u����e����B��Q������(�v��F�WCl#��c��@"3�>��B�pcKlH�Ɣ,�NF����vÈ�JU���*��l�ߝ��$�-�˓[��p%s�'݀�o��|P%�8�� O�M��pVn'���D��}3_���ˊO(-Ht�~"Lb*��9��<o V�@�M�`�A�����A��L�8wɲ]���g*�Vs�� �L�`��}m_y��<Mq%��k�}7d_�ID:0%�K6�0j���G�u� ʧ�z������C7R���v�F	�_��K	���aZ*qT�5n���_N��-���<�� ����4LQ��r�,��_��M
�Ȭw�=0�qs%����_W��q5�I2x��p��ŵ�xV��ި���A1��1��`
o���RA}�/$���
oa�!�I8D��I��^T����F���T�����I=x0�bsF��Xr�/��Qy����R��ǧiJ�@F,1|/�J�B?�䗶��%��x�Ѥ����T���d�k����_�"r�*�o��q��?-
��-oZC{G�95��z��i��o�#�=|=V��CG��kY{v�C۾i�B�|kÁ�, �x��6(�R�
3���XS{��X�rw\�S\gƛA��D����M�}���6�������ε���Iߙ&Y�j�����)]/����N:Ǻ�L�����P������>+�F�DM����籹BV�Eڂ����9�9�(I�T�@{-�V-����j���/���j���m�M"������Lns}� E|s��i���R�I�Rd7�1�|T:%}�h_����<��Q��l������}��@cU��p�-�z8�p����u�}6�%b�q^��f��U�p�w>^<���w�Ke%��r�>�s��bE���Iܹ�A�t���������I��I���h��JdjZ�6�%c�FT�-y�C�w����� �YR�K'�����$U�xd�bI3!
�|�c�| �M41��SyZ��z��)�꼸���R�w���}� WQ*K�_˿\���$F����DqCR�i�vG��	!aӨu�����	p��Ȃ���G���T1`Ȅ�bO(#�$�v0a������dE�!�)(�54�7����FFeH�q�����¥%����J�+?@a�S�@o��Z��YxP�i��(����<��18���X����>upW��$���U%>�$ S֠�ËmN��{��̺�a#�):��ƅ��� �r@)��4����N�s`�����{k���K|��Z�@�]�)='ϊ��s��%��C/&����98����'�n[�����1���Ņ6��4��=������LL	��8��V���Cg�É��K�c���m�P����Q.��t�J�����hz��<l���;R0�2kl�#���������#
~�2b����l�^#���('!���?솄��J�t�,хXlxVHYEB    cedf    1ce0��j�C����t"K�;c��~*z����"��� ;�2�������ھ�w�ϧ�9Z2�]��If�_�$�>�j�v�UK-�;��UKH�Q�
�DJZ�~2i��ط��I3�J,�A����F�1]J�a�ἦ�O�w�(�{=!<�`'p����]wZa�5�w&A����y�mD��;�&�"��߷.r��#0�ʥ0��:e���9"5�!���1�[=�Er^җ�"���-��A=��k~}�g���E-}-b`⽛L�|��^d��v+��taC�do��$���϶�ѻ��^�
����7k��_�V����>��ZO��ɞ�K$�����.7vB蹰K�cE�T�; �g=�������e�z0VW�BC�՞�0s�r�0>�y&?)�,剒�������b6w_ߗ�<޽t�$u�����S�qo!�P�g?R�n��wh�7��iM�.i�S�B�NJ�6:Bf�M�s��W]~�ʱ��fk"�*{2æz\�P��,+W�a:�����b�2���h�nf_`����Z��Sx�B�!���}Mb&9���|�>��y�ޜ(؃!}�?\U�@l�VHb�4շ�r��b����5"\u��	�_�ycfR%���`���`*�:�)Q�Pn
;�XxNC�c7�o݇�囎tE}��Ȑ4tu9
�q��٦���,w���s(���q�hD������#���IZ���N �<�g�/B�����+R��~<MzV7�CfZ3�Oa�0yw`tr��8]V��Z|��D/�>,�܀��>�J�L�2}I!L����u
̙�[�:~"���_V�ś�mIm�C����%�f��'�ԏ~;��3P-6f�Bf���S�(���C.K���qZ��\�����)����;����asx��ew���W?YF���h�L�g��A.��CoJ�z:ȇBc�-�0���# i����a�.�U}¬���å�-q�:�\��h/᧱�4���wW, s�Vm���4!��`ؤ�o97�W`�6�'�w��Ӄ���gG���[:p��S��-5�`�b8F�j���%W��3��p<���^���r�o� �A���S'�8u�ݨ�ƛEq���6�j��6����\��b��.�TșB�У�S5��[yƲ0v'�X�����������%&R��/dN���Oe�q�wɞ�W��(�A����b���/l�"���lEc���/��� �0�6܃텫�ߟ3u�g���P�����#���q�L������O��ᎆ�����R�� m�
�[%���v��U%�a��:�|cq�煻��<��������KG������U�CǕ��dv�9�j�V��c�u�9�O$#VS�񟁿[3��/E���Ӧeu��fS�)D��O�]�����']E�R�4	xPҚR��,�r�)��ʌ]�5O~`U-���T��\�˰�+��m�5(�t��T*
�;���
r͝{�A<U����|�vj^Hk���'r��zj�<h�ɫ!�72�u��Ls~�Q���dG���g�	_C�67�Ő�$'���|Ʀ�x]�Ufm/&s��ɬ���,Lݷ-�RX)�Z|צf�)���7���P���rv��BQ�CуDD��I�=�B����k�٭}rճ�N���͔�-�<�&�
���ƎD����8v�n]�q��6׌�c⼩�z���F� ���w�>�g��}YYW���˖p�纂��1������|x����/c�i��]l��%�6�4�qq��FA��zC���'P1_X�Lk쳾��E�<�o��a;�9;��*'H�zF.Q���1U�^�w30�RVvwO��Y���y�0!�I���t3�ž�ӕ�1�l�>��`W���M}�o�G}heѨ�T����V6J!ʳJ=�.�v!Ff�w^Ʌ
�=����'q뛆|`4�Nl�4]wY�D��!����ݣ~����ݺ�$���9Kt�ag�E��$(��2�S�������k/L����?��w�
��R{R�c5���&�Y�mH99��ȵ��rg۬-� h�uoe�V�@&��S�J��(��o9SV!I	�4���d��4�ק�\��92�>)ۥ�jh���Y	�DiO��ͻ�I[�,�2Wh!ּ���5Y�r�����V��ZL�W&�1b����Q&���[
�/o�g��$���V���W�����6	�l�I�2Qq��n�̓����u��k�/c���
����uX�h��|��؃���
�3�D5�'�Ӎܨ%6��&�ލr;�OBy;�6�F)����� �����u���=����+{ʱ�G�'��V�&R��n.��ص(�iS��<�V:)�����n1-�����]t"��ⸯ`������T����	�
��n�hRR���R+�6#�8'�&c�u���T�bѿ��Q[흛�Hq0�SH��E�1^�.�[� HM��^�#W�� ����
@��O���Z!D��ޅYgN��.�����l�b���p�� B<��P�fڌ�=cx���lʿz����Ȧ��B�n�h��Q��E������ԋ���g�&�AJ��*'Ƭ��='��a��qj&l���i5o�Jp��
�I�잼#�%�m��yUv��1p		rN�B蜨��!B�Qk�~9���I�.�EM�"!��Ylv�*�����<��k�i�#=��5C�SkJ�$�,C �ϯNa���xi���as�w�n�/�2�yc8S��7Ф>�ʵ(HaV�E��=W�ɞl��j'_9	��A�7��c�G����>*r��(|�o���T�[q�laI�@;	a*^���O�*K5Ž�m-)X\R��e�M�ɒ��S�	3_K5'Z4u�c��g�_,q�w��b����b�A�O�؋R�Pu�I���\��ɂM]0�W���C/�h�?'fu��ipʙo���u{-(�o��t ���\��':���ޝ�j��]�x�j �\�;��-D�*\$�Y�;<��o���;]�[�K�v��s���O#>�-�(򒫇{DKA9��G֠�U�n��������^R�}����Zx��{m$A7���D�d�Hn;k�$���{O�t$�gv�w����"�׭��.��r�]%K.���/��?�/��[ϐkaٜ+;`��g��5�EZv+j�>�A��R��G�LvbmP})y�`҃��ʃ�� +�xo�R��Zi��wz��j(]�+,�T:���? _����|�Y�J%���~�q���3�\���.�kJ��-c�)◊l[���f��y��WK�5G.����4`��izD�Ѧ�;	�>@�&gF<c���kʏ+��C�9��/������͋�x�dCץ����wP�ְ�H�ZO���2�|7E���k�1��t�0��D�s�~"�Y��!Ot��@��!��$�+[���y�8ΐ6���F�E�7�١����	�U��}]3A|�gTOKM���?U�uرK�@\ Q$Qw{ Z��.?��;��.�ףFɘP��n�m��?յN���&n�I�[kvu�Y�
>�K!����+"�U��^f�-j�K_�� t� P��w�d@Q$��m���y���m�?\��L����&:w,�EO]崁�m;ccQ�EQK��mwx�U	�w=_M���ɽ0a��O�s���+^Zm
&��+��'iC���g�=v������%l�0�M�oƝ��'nQ)�?��1q� �¤1 ��H<�21�����0!���/^��ON�k�?΋�� ǟ�x}A��8	u��l�3���o��W��;���<{k/5$�~�-��,$1�g���u�zx��H�����5	�~���Ý Ia�#�x�ٿK���G�i'%ſޝdZ��C`̰��h��l8#.㻦0�cJh~�
���aV$��g���	��?WS��͎3�L���N�lX��O���e��^$�R����yrd��G�4�M4c�+�3��8�ڨ���:���^���_D������t����HD NU�L�P�_e��lh����72B(��UU�"��ŗm�S{����1��/��&�jzmjس��1���K
�1�V\5h_|*~�#���}OUA�Dô��W�]��( b���!�gS��_`�o��Q�_�3_����t�����K�˄�
<`a9���5�x�cl&;��b���oGQ�_zm�_gZ�f�
�,�+��d���y���&)㑌��+��9tZՙDi��b�\���Y�������\�Jq
�x{Y��%��8(���OCɘQ���5��H��^��nd~��P�[���Buצ����-�֕nd�ȭLP9E�a��e�5m�#ǙX� V뙮����2c��_80�y��b���\��or�Bw�e<$^NN�PM?���� \Y���/bPu�dH��<S9��}βfO�$�-kb{,�:2.�=ٺ����:p$�]0?��=�_	����v����x�@���ď���o�>�L����se�����B����"�<���&�t�t�Q��(N�j��TB:|��6�$���C�.�_QU����6��ӥ�[��X��1� �p�M܅3���!�d��������x:%₨�����,߆�x#��&/�J����vG6���A
F���`R0Ζd �z��/?Y�4��f�x��Ob暴k/�J��Y{�tVD���K�ȵ7{2c�Ã3 �C_�j����σ�al�����@~:�Q�7:�$��x���^���g�m�T䉈�r��&&2���T�����I��is�Um�'Q�"�i$��tD�Ƞw]O��>����R��P�~@�y�F��2I	j�*v����j����<�T�Ӌ���S�ȋQ{��BSu$߽Ūۢ��B����~1H��ݭBz+�ώ�(��P��h�*��XZ�@��1�0���yO�6�K%�6�0���������=�GA'��#��e�TTC'0��Hkj����=1v�9AM+YT
�,.� ���1f�Q�k��ʣ7�X6��R�|	h��g�$�-΅���?��e��8���3��A;Q�<ݰ ���8�l�L���?��RKإ=g�sÕ߇vM�����&�gs����:��v<e��+�G6���'�/k��=���3��2��j�{�7��q��R��~�B?�H܈��=p����H���b`v[0�g��e��o?�Ќ����:�iqa��J�%zjIq�`�b����&��^�����qr��u�<zK�F�D�Fw��|�@x1�B�a�}�\�T�Zq��)a���2�.ɉ�T��f���?}H0u�v��΅��n�=�p�N�9u�y���. �`8�m�Ba�W�#
��HL��ɂ�pڄ�^{��Z�v	ݜCc�-�?��\�t��B[˽~4P�i�%/�mܔ"�u�aX9�V���S��ٔ���<a�I����Ͱ�I�zIN��X���Ƚ+'g��'ʍ��d^��`�ɣ5:�}]����h,:����]�w��n�Q��#����K�hp^큹dϏ�tFz6ƗEU6��Ӫ�rV�~�S&�s�6��HR�~�����=�nJ�_ɚ%����*�����_zL�4g `(�M��R��P�4Y�J��-���#�o\�|�ui�0_�d�q�D"ֹ`q��H:Vu�)ۑm���wj�-��x=�@�IRG ���b��Ş�uoz:/PI��B��?3G�:�(K���*�"4�������#�)�k��`���7�"
+��!�e�&�7F���m�h�uEc�{����6 m����pUW_6�|�ɲce�����]�7�
�EG�l>m ��u�[=( L 1��p*Ɋ�<�8�ll)z��r[�^?��qg2�˟X��KMo3j������CQ�V�#��fh�)�7Bx�g���.䩾�Zp��,�=ɱ;��Q*��"V���)�'�MM��iz���s�g�>� �m/:�R�I`����^�i� Ԭ�����*j؍g����~;�����6��G�xS+y�"����r���@���&�6���?�TE�ك��H�ل:w��E6�����Xû��e_pz��;�>�ނ�&��L�핱n��
^�cd�%6�]���r�`}�PE��Q����L�,���G���2��i�����(��Q8���Jӹ�"b�'3�D��h�:-Pr5�o���E�����e�ugE]�~��9�<s��xE:+�w���y��نP���|�ɻQ��'�v۬z�M��-]Uu�#�����o����)�ؚ�B0��:WD����,'�Xp�xW�`��l�`�#�5��:Ňz�u�66 ��a���N�->������a%0��;IK�s���;y��DSl���i��7J�?E﫛��_�J����O4,��/v^ !�i��)g��?��b%�ٯ"�Q1,i��owh��+�(�k2���!~���b����~�X�?�kq3�F���+2��ƞp^�7@Ǩ�zN�βBg�~[�js��_1N4��xn�w�1�Pn�#�2��.6�385|��a���+�����\���u�Ζ0�g�C����\A��'��𪚮�>���|�Q���Å�d���5=�n7�Q���f��w��mN �s���ur�T���V���� �F~�2%���% ��Px"3Un�����,Xs��1N�_]��ap'�I���H�݇İ?�/*�F�cv�. �w}dԡnS�ۻ7��L28�ĝ�]��.ƪ������P����V�8vDr�fp�d����ԭ�{�1k�ޓ#w=h-~��U�s'��<�;�gmMB��B�UuX=��]���!Ds�:B�o��RѸHϾ^��e�k��`��C��DHʪ��'_��L�b�û��]���E��[9LGR&����Q�u�aV���[:��x�s�m��2ߺ��ȃ.�_��i��po;�)�=�j�اF���t��&�>�e	3c�2����}�v������(���=���/��_�z�u9RU�;�ʀ4��4
w�`a���#2S���	s�U@��ɔN�<+�9�0Պ�&���ȹ@��w�ቆ�;d�5�`�����+�U�uG�4fv}	�k������������U�xj��s�G��ù�Ud���S��-�޽�!v���H�IG+=�qۢ��26x}?�����g%x7��RB��^�}1����f�F���ԥ�A�ӔY0���(�