XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E1}�9_�:#�ƌJ�ͼ��� BǢ�K҇��M�p��>fB��ݥ��)ʦA�B�Ҁ�JmK<���)`o��Z���؍���/w����l��l�S��Rb�\B�o�Nx3��C��Q"�� ��v�~i�<�����L��r;�ƙWR���0�m]�42��NL��DLMJ�7>τ��hY����'�[�+��[k~�l�)r���h��u���{Oʬ�,�K�|���3����B�X��;��OyB�xkcK����� ^"k��uI�^�9�ӥ%~��^�l���f[��\�-&�x��;��R$�e�Z2hD�9���d=����m�E��:�f`Kӫ�>�O�Js�(�6&�8rKTU�y �?�"=,to�~�[|@��¼�<XKZ	&�7m`�_W~"�ȿ�a��K��[���]�� �&Y�#_U)��� ��%:yM��"kHS}-X��JP��;��:��`�ArU����ɽz5�7�D}!����z����L& �̞�1�\ٚ�8C��L����yy����������cU(:��	�V���#!QXS�
W:����ڲ %j�e*L�(�vZm�R^�`���tɶ�{)��7�\>Z�P��\oE��m�5����/���Lk�[yD�oSwz�mW�O�19?|,��o3Ь�.����;
6�l� Dg�:l�����r{%r��9�/,��a�%�����w�e� �iJp"ae���_�\ښ)ikNꑛ�7lK-XlxVHYEB    2042     880U�լ��#9�����l-��Y.�ӲIR&�x��a�Ɗ$���\��O��`Sjô���6c�"�kt��x��1����&�T���`>��������Q����:N-����Qϩ96�Ȭ�Zq����w�_c|�g�Ӕ�^�k�К� -��pwTb{zL��+R��8��"P�����[��ecܽSpK��)��~�Ӱ�>�2@�� >�vG�	������0)���.�xA���Csy�s�H��_*t��ɀM�9�}��Ӊ`۲6PH5�57�`QPA���b��F͡�@�H���؋sգ���ׄ�s����/��=�jZ���o�~���;_lD�����s�X��|�Q�HC}���*L�Il��59�0Zk!����B�I�8<yr�t������H��ݛ�m`����*$��q��
��O�%1]Wmٴ�I�=q5SS����&n�a�ۻ{���M޻V1�g�Î[fd�c�e,9�:�xc�叡L;G��Pl�.�/\�!\�ۼes����������|a:7���7�`��\��TĸR���|��������;x��NXgska�9qKR�/�s$�U��Q���ʍ�T�����g����4���?2ta�SQ �*'$�-��Ț`O@K�<�V\@�Խ��� �J`*���۵e�Ɔ���UȖq��+�ETЏ6W��|��bl��*�	�Cj�K}�3 ���0/\�5׻xF��e'�.+��ZVҏ{I^��S1��;�ݽtOs�U�������W@S08ZM0!z:>l�� ���e?o �4ݫrM�G�ܿ��v0֪�dV��\%�q?�n;�l�]�B� �%���oPD����k?���
��H��~X��5Í�����8an%��n���gC��2��<���������᪩�0�-�*�y`ӟz�^׾��܆���g�ꩊl�����Q��e�f�{��d�p��K�l&c/�qL��L/��t���ǭ#YmQL�<���zy�N��d�*mݤ:2.�W�T�V�m� �ǜE��Wa���n�z��za�� RZ�!?��n`OtG����)��p���ϑ��z�Y3�TT0?%��������~Fuvp�[��$�"�xRS7�37!c�n;�v�Ն�܈�� E�ʓ%9��nւ2v��ٯ
���E[ߜ]I����-�'��D
��D+c@*��c��|�C�@��!�S������e� ��KC_�9���ݨ$��&���@�!��^�v�ؘ ����؞�s��4GA_�Ic4oZ7�9g��̂�U��[j�BZ������芞�_~��Ջ	Xt���(�\KP���a/�?k�>)�z���I{���"3CH�s����\����N�B�Z4ܡ�����(Z����!f���z<$��9	/B�Mh5��#x.#�h��E��#guT~'��tA�Jo�Öuc��8|[g��fV�|��� �Wd�;���/p��T<U8xթ�i���3 $e�8��A^\������B����]�5Ci$b�0�ӌ�9��Ea�2��Z��G�A���N�cJ��,�x���*�	j��Z�c�r�5�
�Rz�7,R��a$ǳH>�s��)I��m,h͏��,FR!i��N��j�Ӌ4]�$�D� �s2�� ��M��<��N}��୭)m��d����[ih�H'�X�,e��qu�O�������1�δ,�*$�şb]��U�xA�����D�R�,�yR�B+2H�����z9�M�.�����z@���/������Gt?뮽�p�3�L�tz+:�-��k.M��Wx��]�)`.��qZs3�i�J�\|܉|L��l� Uo3��>,��q3hpcT451����	�7u�tGΊ�&��v��S4Jw��*-Y���>��x�[%3fa�9��a	�w:��İ_�+����^�3�]�l�h��9�@7��l8V$/��}U��QR]�W�>e�j��a�$��x_U����6��/���c�^Ԁv�3$��Cd�	!񞵋��[H�(D����$ل
`?�w���X��ٕr�H��K�?������j�Ǔ	(����7ޝa��T��0OX�E�N��Z����( 