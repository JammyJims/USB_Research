XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F�����dAj6�X�����{��/�p$;��-�_\kQ�z�O�A�P�@�<wP]|\�,9�ž�{H���9UP�|B͒��\ຮ&Ƞ"a裨�a\��f9�ts�Oو.�ʔ��kl���0�߾���r�m�<uoZ~�����[`XmUy� !�W���S�B�o�dE��sPz*��� ��+C��!�xs��ȅ�S�ʖP�{��ҥ��AHUbAtzD��
�#��)l��9�M���m��g�LT,R̔��6����Ab8LAY�>y��a�pXD o���\`)�5�VĄ�f�����6�O<�W.uF��0�j�GR�,;�\���n�,dR���ü�)��j<@���ƍmC���꣸qu�+���Mf�ޥ���%������hi�r$|�b��K�]�Z�l�E�-���x�*mϨ+ܘV)/���z�� �?��;׷��ʨ��Y���k؄M`,��Tv3�[��8LZ7�L��(zYO�r�o��kX_�d�a�%`ъ���S��rL%`�ˬ�BȪ
o��Ӱ߳ԍ�5>�iTl�!�>���f���
mq�&f��`0��Շ1��
�&��բ��2���.����=�����H2�\�>����9��k�:6�Ɩ�r���x��Im�t��;�n��0�RIS�(['k]a$7�w�@�Ɠw�uVRxr䞊I/�nĺ��FWv�"Ų^�8�(F��,a9B	?�zw!:;���cڝj�!��f��vE�~ՎXlxVHYEB    11b6     740��l�g�^"��9r%$")Q�I��4!�ыW[ЇL�^�����LV�h	�6 $I��.[�Mg�9��Q�����gG� ��S]��̙���HȊM��~hA�Z�/�	.S_�����Ǉ��ź+á��G�N;k͎n�),����	�/5zp�=����ކ:?���IXKC�j?�y�	�S-���� ��2�0���]�/D���{���.yGUC���Gyb�r�MA$�^g��ǖ0Dn��*���Fj��i/�-��*7�&�_k�� W�>�mS��7T������CȬt�}�l�ҥ+�f.�^�q����#��y���Wص�ij�*y}�蟷�혘�s�A�*���Md�.�@ja,+lOg�� vBd�k�������G�c���G������y��6^�x�6V��z�?Ւ�9�U�z�>�;N�� ��.@[դA:�A���t?�>;Ԡ���P�e��+;�?2~�$�S�EJ2'����)�16�?��d�~�3�~�+ ��b�;O(?Z��T��i4XJ�&�%��/r��'?/�Tx-OBr] ����kk)�WF��T�N���]g}�%����A�e���)ʃ��[����,�]�,X:JŐ�l}�>�f���7���֫��o�{��q�UXX�;�f��7C�ؑ@'Y�*���y�r2�b��w��U����.��I��P�����Pa�C[�dP>I��;m���U��1o��E=���6��<��q���'��hg����s$��ܞN�N�=t��S,c����/�yt�$ƽk#_����o9��ϩR��}3��;�\Ux9���ag�a�Z��ɿ�$%0��T�/���bB�������Y�PL���s�"��
�~�����ϮO8ԙ_��u��#���j�o]�k�ʙ�A�9��b�	���h��vo�Ex��RO�CQ(:򮼭�{���/��'U�����+.� @cP���p�&'�dM̘@m������v�0O��F�fc�_K��S�H/��߭�oo�#l�VpN׬T,� �<��a˿A�'?�|@��I.� ��Fr{���N�������\��^��S�0BX�Ƃ�Ǚ�D�1�v�l<�})V��s`�9����O�Nf�(x���Z��K�W�O���Ǯ{o'��b"1/q�,�/a���
��W�e��H�} �Mu�):(P���M1Vj
\��)����s�[�o|&QP�x.zMF��O�=�V`�k����7�=Mө!�}h�.������ye��cJ2?�m�U=\_Y��t�J��݂FeL��� ��l]�Lc0 �(��'-0M��~�B�ǿך�7փtt���+��e	��Oy�؊[1G�Уs��H��5���,:�4���"����$_>�Z��u}��r���'��
�h�)kTpe�?�Zgz���A��ۜ�qp%ysb]ą�G(��C$�r��-�1q� �v�옷!������%�Y�p󧔏�x��|Ue.P���� 
����㎴��x's2��Vd�g��`��Osm.}��t������i�&��
1�B�r�t��*A��>2>��W����l���H�آ 
����V�7�?Gš6>��θ�'����;Q1E��)u�H���#���Tq��FF�mԷ�>b��;���39�$E��jz�R��iP� A��B�d )����ϒ�����+�w+&׳��f�"`CC��I3���մ����oDI(`Sg_-���~��/dʲ���µ���B��&N��̮'Κ&���K�qT)f�=/cx���