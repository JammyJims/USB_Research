XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{����џK�F��O��Bo�n�O�;o7hC`Bkx��CB�M"�N�୧Ž>Edվ��A�?��2`��+0�H9�<�4-�Pk�Is����Yh�kC��bѩ��N���ʟ��Z��̝�L؆�k�s�Q����Ԉ#��z�
�76U�Ķ�ؠ�����$X__�f��c��W�0�@z����}Puo8���"<F���ޫ�KW�幑3Ti�>[X� e�޺C]-ϻY��z#�������~�.{����z�쁧y��w���ҩ��z��@ � ��j5�?A�wK���RN_~W��2��8�����3xsn�_���J-+�D�!_�X�P���$��X���9,�D�>�5�x	��V��T�tv�|�ʇs�{�(�ï50+B�ɮg���u<_^dM����BB<�=k}���� i¿���d�e��"rv����i �\�jp�Ъ�=�еXi�zY\�{��.vt�	R���r�s��4Z��I�9Pڃ���;��$����z�{Ы��x��mA��D�����Ypo���{<���=،�=ÿ�6��MɞΥ��m����+�H�r:mawv��y֎'x�W3������}5wg�� �iu1{���x�(�YMD����Yj���!����r�3���li�&˷����|%��b���3��j��-�S\ �|_@���1bZ�a8Md��-�A��Yd���6���{}������W�_��_�u�6�@���mw��XlxVHYEB    ed45    24c0�pU��-��G��V�'p���U+��\�!me����b!14��$/���ގ�3)�[䉅8�"sŎ�:��0?8�_���Ψo���jI�]��Kf�n����Y2:�r6�8�e$����DU鿬���Y�[�$�8�6>9�$Jo���=�𻖥�Ւ��߬��|Ezs�!(���t,ר�	��y��_C0��w�x�
�!��p��PO�|��ۡy� �I�/���|�v�s6��g������ |W���+�w|Bh�w�-�y\��!�8�I6t F�emxD�[�J@>��Q�Y��큕_�~�-�B�E13J�t~�>ɍ
���0B���2R �U����_=���>���|TT}��}�y�O�2�����BW�~Vf/�: �-q-8SAw���A���v��@�$ͧi!�)@6,_����؏#f�y�߰�$05!��_D+f�c��8`,h�a�nt�h"�F*�S}b��A�r=ޱF*��j~����8�9I�wC�b����
���i%ƙok�d��� _�g��F�0�ni(A-��ot@�C�JY1���]��_f�Aۏ]+Ol!�%�u��"�Y���^��c˨J��}ڹ�{0c*ݒ;l[����C�d�)n�2��^u�I������<�\b�UQ���p��"2߲���^U6�������Ƒ�Bf����������b�6��7x��VKH���g]N"{���Z w��g�{��Ց19C�6��U���h�>x�[[�Hӫ�V����De۾�_��UIo����ZD�>��y��]Wz3=%�PH�%���~ff�A��>m�QC�w����qw����hVc��+�_������	���I4K�"H�oUvG:S�e.H$��3b�h/�}��u�j�$�׋Q�*����5��|���0��b���9����xeiN^	iO_�[J�����b}���dnK���}�
�p��%���فI��±�Dgf~R����7<gv��%�p)���G�-�+[�(���(�9��P%~��Y�B�W�F9s*�i`�q��iO?��b./��i�N���li�{Kʳ�I`���> +�/�7�/����7�0۟2�?�X��0�r2ڝW�"�c��I�fU����0Q�V��`'B������CO$hi H�3�/�Q�J�݄��\6�kkو����8�j��� ]!�q+l�env��Vn~�>�w��e�>�rĬF��І�8�Ԟ%a��R4 ����=���_�24:1)�:A�uۂ6�[��dk)7K�a����o��bl��af�������1��s]�6�ZXA����^Hٓ'XV�N'?-p ����]�*p��A��ō$2�IHՋ|;$�,�I��H��<�Ҕ�h��(�f|��M2P�hÍE�Ϋlߨ��ıL���i������G��]�?�A�9�m�$L�dNn�I.i�I�D$̋Ձ)3�a+�r��C�(���/�Y� uRm�W���8�D�[��;���u����Cm�紨�/p��ht�:�EM?V����V�ޱ�����/��-cD��眾|�^�jC�,�.������r*�	��D����+:�|�'����K�V�R��f{n�Ze�Z��k�)��ú�
7��ɖ|1�ڤb�T�)n�1dj2c��?Q��(}��yzK_����LSY���BW]#ۘY´D*z�����2:&^�4q8��_��D�k+ۜ��:���)��^�}�e(|�IC���3ƨ���8���*L�`a�d5Р\��NIB�����յʀH���~�X�����F{/�1p;���I�va�@�AD�p��wO�y}������l�t��UF������4�w,nm�vҽ���u��^s^���;F�y�i3,�"��E��wQ�0�8vbx9�O~ �a��	��k�r�M��?%��|�1�:�U1C˝�,����'���?�)G6����+buCW˄a(^��9�}�W��R1����}MZ�ș�?��	)��Xɶڐ\L���ew
��K����ŵy��"�Qӎ��z�$�����O�"�|�'
/2]�i;�O�)��������,_!��b�5>ѸD������P���R|�9�%��Y'~���){�",ȱ3L��DY���̥<p�mg���Fμ>jrѴ����H�_0A�.�[���<��F�'!��b}Q���"^��y1�ؽO�l�/�"|j-v#��>-� !��v�>����8ِٰ����l��b]r��TUGQ-�h	�?~� f��I8c ,��1?�czDL������"'Y�"5�8V_�A��S�4a��#�29q<�Y���wXe��F#3��9�-��w�1o���bB��\~p�׷_�#TD���1���W;y������ڮS�5�xQHK���YհI5w&���:�ĽqӬ��_��L�
���URQ_�/܁��t!����;���x�d�v�m;
Qpϕ���T_�٧f�&�� 	�B�+�C}� �v�_�G:S�F�A�=���t���o �Ƀ�MM���]�������+r<$C���r�+Dɠ�gS�W����R�rϿ�*J�����T�ʏ��JEs����d-'��(�غ��|84k�MVa�W�Ɋ�B�}�G0��?۞��e���z:*sEO��Ҽ�������D�;��Q���J��"�@��"���q߽�A�1��"��X�ز�����7��W����xٙ��9����Ҕ��{��<�"3Ia���? ��ld";hDPf潖�r/e��d�X�R�?9�����11��/Ew,6�O[���ב�M~�/+?J؊94X�!La�D��<Y��'4��8���i��3"P_��'��,���ٶ1V�p
Ǎ���2��3�ƺ}��}gWM wb��A�Q|�Z�֚��~��� `��Kdwqѽ�t�¤9�bb��[�#�Q�c��(�1{�����x�:Wx!�BAIQ=����5F�8��V)��_kB�|��׈rGԑo�z ��^hz�A��y5��h{1U���_�O��a��9�����Ž˛�t����W���H���<0��%Dtڊ�#xػ��OU�$�]eb��G[�1��8C0�ӝ��<I�9��n[W
�/OS�hOK����Dҙ=�l����V͟���э�Q0s�J��Eg����4)�[�!�Jz��j�`��զ�!�2����V�]���|K�5��54$�S�>�{fe㲖.B �����ĬX�A|��,���̗�l	![_i&����z��ft�(M�+W��H2�#$�]#c��v��MWT��XU��6�?�B�
�LMF�3�e=���W:\�~� �x�ۿO�jk�J�4��nV��S��:�~y1��(�d��q�����+�����[�!���g�A�����吟
E{*䔒��
���m,=�T�A?��ar�G/�]�T����I-���\V�����ӕ~��9�7��wB&iĕ��қ��Ě�$�+�>�׻��q��7�a��{㦡ѷҬ�O�B��tմ��p:1EH%]�a�0G�|�IU7���O�Ym5�:�P�#��ں���t]�����"4 �*@H�F��yx6�A��\�b���5�;��5 ��@�^)��U`G*�û �L?
ż���.h�ۗ��937x k��w�[��ԶNl�KW����<�U=���h>e�ҡ�ːtR��� .�v�?{�k�-�yUF%����,�r[������0 �tv��?z\/� �L��l\��.fQ:����/�,��Z�]�V��:A{Nu����
M��l��v��)���Z(�Ⱦ�~dP�X����_�QP�zPi��<�h:��hOK�+��y.|��[`4���>Bo�~|Kx�A]�OU9�,��D���e�ͻ��B�Q�O�x��
N� ߶�ƺ�������䛾Yցo��I�ْ]80���i��UC� �6���~l�"۟������ù�QP$���G�2s  �8�cJA�?0�2F��E`�)���p���z�fU{AP���Z����E���)��A�C�҇y��V�����\%�Ky,�m�%��x�&!Y)����5�b-Ǎ8�r_�p7���Xݡ�P���,���6kU�=�ê��lįDϘ�sL�����IV��Qm�y~7[	/���vӶ�I��N2��'����� ���O��ZU��K�P@��t��w�7���Xs�a�?^��#��ܙ�ɟ��Á�6�(�P@�{$�����V�������B��N'�uq.���׼����Er��>�ۺ.{������0��&�v&JK��N��XB)]��g�5�W����fר���#0/�E�P؆�Z(c�C�p���V.r�vc�Ah�"�o��$���H�~4�����hj5꿜�� �p�e�'�@����>��99���ZP�I��:�(��0 �p��W�;P��`d^HF�_1�2�dk�zYo����F�F;(�Di��f-�	LV��C���ݓ�7a|[���&-�z+od�#�h��5�^O��8�~��)6�VN��Yh�R�v�QbXb|}S����?N��D�7�������f��k�Qj�Ă�����=�}�%�Sw���r��(n�[9�c �'�rމ���v]�lѶ��1t\堥ƘJ����Q=Kd�Wʱ��ci[U	ޢ_�g���+7OM��%��a��jx6)*>$���K4��5���=&������`4�r]�0�f��e�7@�R��վղ�(����z��e�8[$ �ʸ׀L$���	�p���=����07~�H���_ah�O?�v����Bi�B�n|sm�,�G ��v�OX�/����p�T��/ѻ��̍��^��^�.�e��*��b��vZ�O��%���lj��Uk%�K���]�r��t�GA%���ȯj��T|T/}o���{L�P�̯*ٖ���Yyѡ�g�/�� ��t5�tϚ���@_{�P�kTC�J�٫��G&�����,�[��w��#H���]����a���N�:�[D����ͮ��m=�A]�!	�#�̴��N�*IY<�P�p��]���š4<(�K��^��pC��Л�H�gl'�h�~�
���nǛӋw�J͍gP3I���(~4k�-#�CN��ze¤qZ�,"�m�HД3�@���ӛ ��o�vۈTZh�;��z������n�.�u�x� ;h���&I'<s2��y��K���IMf,|3@�.�"��G� ��8��2�ڕ����q�a޲i��i�_~p� i׃�Ӄ�)��6
C�v�HhY���"�����-��)d#�����J�	j��`Y�c�ɱ���{�*Pc��za�	u�H+�	����cg�/�ҎX��L�뒤�|,^�6f��v��@��>��g��Q%aV$|�!܉M�1���8����^
@�Q�b���X�۸��D��*?y�<�������wh}�3��F�y���_8��XA[c�_tAZ�.	�|zx�8߬�A�l�������%��Nj��J��)��g�E Dz�Hzi��ʂ��4I�a�M���q[àUln,���7�W��f���C>d�׶��"G�Y~u��q�X쥜����:��WS�^�&	7>����pJ$��1�0��T�\�]��M��](VsK��a��x&�֭�DXf֚3�?����mQ���vn_�ޱ\�����o;�� /f1;��}y�bK!��� Gr�= �V]&(���=[�u1�fc8̫G�q���zj�$b������K���9��&��"�a�pbCb�3�4Z��a��\u�<���e�w�zT�^W@kt�U������lǐ�y��p };A5ωFw�g��Ԙd�W�6���QnU/�*�So�K	���ls�����2C,�|)GO{k[�0yA.�X�T���l�J�J\�wG�0������/�w�d�#UqGstǏeG&;�\��CxˀxopQ��?����&��cY��{���4����m
8Sq#�s�����U-�R�.V�Z}<��	���I/p����J�C��{dn��IyX�k�Z{Ո+R����5�.���4��C.��}���Q��0�sh` 5�|Yx�-L�p�K�{������Yw.�~Z�k�=�u&m8u5��O��@���;��j�Lk��XX�<6ሉo;��'>���RJ7.�D���8���3�Q��A9��DF��#��o����f<hkbp��\A#�y�O�IJ��]�(t�u�*ڨ +�(�gmt�e w�y�{A� b���h���$P�dx�x��ގ���m����o���ƿ�d��R��l���{mTCz'��\�Q�X��P�I}�~ �.wx�����(_v�c\�Pbo��H���cA�T��(���תޙo�W���g��P'і ST�v��g���q%�8�enOI�r<>	A�@�>�ݛ���p���=_�Qr��aI�[\x&��[+� �-��g@�y���6�ƻPi�,lu����z�_}�p��Z��U�����_h�O����F�no�Z �j�"��P���y0�	J�g@q�j<Fǡ͆P1��T��@A������Sό����ӓ�}><�3Y���vU��q�]�2�n�F^uɫ�ۻl'�>���S�G�!��G�.Z+scpmֹ�w9>-K_�2<O���S�n���(��,QO�w�T\�5��ͦ�2��	)�N^����ۢ�2���@�-��.��ǉ72M�������Ҳ�-�e��ZܥY�<x�w�3���Qx֑������7����=��XM�4	���D�SV� �o�O�B��_����3E�Aܳ��G�x4��W2����ӆg��"�k�mP��;���Cy����U#��ʐm���O:�a���^����5�n@���/1DY�e���5d�� l��� �{��]�!�C#�ˇ淆F����9����@�`���[J�yRw�=�%g#����˶�>�癔{��S�m{k��x��-�-���}��G���W*�5�QN�A�@F?V�:��֢����3_~(��R�^�[��ݛ�̳��<�@����}r�P���k�`�#;$+CiTk�L����}��ʹ��d������о��*�8��q]d��Ha�4b�	 �A��	�а�A�nG�t+�qKɽg�4<��Kr"��~��%ۉ�MIG7���q
�?����"A��H���oh�r:����@�4c�� Մm��)/��&_���
��I�(8R񧛜IF�
�IRVzg�X���A^��H�>���I����%���E| m\z"qG�M��z�kXcN%��ĝ�M�hQ���	Z_�Y*^X���g��qjX�r]=xrpa��3�~�
8��rֵ�l��K�[��.(R[���#I��-��m��3L�v_*�k$�� ��=�H+U:CO[E����2M]�����w��w�-v�8蠚��8*rw���3G��[��6��F-��/]x%A��q��2Ǻ���q6Bz�����#���fpg��W���2���� n��~`$����F���17��d;JR}�U:,�^@N0L�u�I��h��&���"cl�y�D�#���{mۯ�ؤF�肪h��}]d��U��a2����̲\ Z��C�F=-���!Ao�v�G�Õ���h���o�K�w�^²� �)58�$� ��>�f`����r�8��W��n���h5'w6m�e��YW6�6�M�ե\o�Z�|a+�o���d��T����F)Ḋ����[.-Y�J��%L)�}`�jV�����b����"������"6P�l�4�`u��FS�Kڢ��f����&��@��-�%d�����6�h��Xﰵ B���l��o{���Ov�-O�R��R,����am�:�ǅX�e�o|���Yڶ�~P��~�|8�|?���%�{�%�U�O�.Q�a@�_Y)}#7��f0�'17���r`���~ѵ	v�:�"t���
"���5�ŷg`�oTF��	{Ei<.�R�-<otulM[�$����y��yC�U+�+��;�-�'�r�F�p"4u�CSh��ж��c���ov.B�[|33���y��	���m/�@6�u'n��E�������xo�0����<%	�]J��{���Q��@y4���\sq��ɇ�=rx��k�Q�7Z� Y]�6��d"Oq���yl�kN7B����p����,h�w��� 쫢yY�߁����o�c��o�K�$,T�x*�����vsZ�����6�N�Qpf�G$�B�Q�BUmА5�gs�R|���W�,�K��Dd��S�Ř&�#��-a��:��{��	�.�ʚ�F3�ͥ$�11��§�'��d����V�qi�g�,�Vw���J��fN���ޒ���XבB��!�L����������eL0 � ��q��|�ܼ1{����~P�Ƃ=�� �&��:X�Ď�����~w��\�x
B�����<���@��Q�i<��h'u	e,9�x�?�<I׽�Q��IU�z�A���>o�� 9�W�0]9q���Մ.V:U*�S�[�v[%٭uj�mE�������d\�\�HZmd�,C������e�#n�Ǜ1���D5�� ��dz�'
�����ҿR&·ۑS<�����w��P���sb����<c-�� 6�8�?��(8[h!i6v�n;������-=Y7�P1��ٺ�C̚�>za�fx�b�U$LI;3	Բ�fB���Cλ�|��=���g�m>�\b���#������R�1��fF�HU�'U�/m�5r�v,�F��a��q^o��<�`�O�ֽ��.t��w���/r�oZے�!g^������+����M�r+��Z^<X���$�xl;��3Y�4a㓥9y'L��@����\�"�[�z
�P�]�JM.�
w��Lb�zԂU;����35���xFQ07R���n��Z���E�����1���ص)udHׇF���D�=(y
�@Q��1�h+�d�3u�,A�6L�
�nF�Zߙ��K�j��ʟRp%���j^.� ��� p�u^�m�t8(��{ƩAA-r:pw~b�	Jm�����������IA7�h[+"N