XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i���k�^�2�#e~?�@���(����F����l�dsu�/s2(�âq��ޏ	�����ѻq���Bb�:�٪(ِs��D����c��(ǻ=*�DF'p���0gI�D�NW�m>��hs�������X�L�S����b�.g�c tv��<�a����xCL���uf�P?�'X���w�6����½Dld����\�!��i{�wI{����M^vvv�{�>���n����C!��{ǉ�����Y7i��[�=U��gJ���<�	fչ���R�W�L�1<��l�VR[�� FxS���#���N�d���<��83�\ao23�s$�3�+l�h�4�D��ʮ���� ���yW�FSd��l�͍�M��Ȋ����W�����]��`�g�4����I����&ϵ��p�q����iʦ��ʐNt_l��S�]!�"����o%�S��6���"�o�ل�ymupE�_z���DPR�{�c��ÉgyQZ9P�e�ϔ��N��-7��I-����he�5�H�N粀g����!.�Q8"ώ��ݶ��5)n2��y�'����,��m;����T�1��[D.�!0 L ����8������:�6����v����q�ϝ��Θ��!�x��Z��3�J��R�o0�l�D���EEj�qC�W�i�"eZ�����M�,9PۋߑyE5�s���:6yP�v�̀��}��r	��(�;��I(rVn��v|��>wXlxVHYEB    3248     f304�N��Q�X���3�����/�+T��e��L�ӿ��j:����1@�uA�v���"'��:�T��\g��`=I]�}j�Wm	�r�Ð +ܐ�5 '�Ŝ ��C%�P�s}~���Z̩!3� r��
S�����Sr��9�qd<�t�.��sаC�� 5k��L-����>�$���}��\r��l�
����?�f����X��)1��?j�Wj�:f܅\��1��4)�F�P�QZX�{q%��okbzc'��v�^�to���?F��B���ֿT�'|�ʴ_b�z�N����]s���eOJiqEC5���*Pmէ��(/x�&��V���huC>�W|��7�ǂ>����~���s���tUR�m/̟lI;H͗s���x���<�~��[�r"�ZRF�g���"Ӿ#N�eF�fi��
�G���N\�(��s�4�J"��3w�"
M���3�)PHt�B�1�+A�j�s+4���h��Fp7���y^�<;�!D���?���	g)H>4�d�wvc>��Z�)QK�����gʜɨz�f�8w�.5�	&ϲ�2y=�;k�+N�j�t*���k�\�3F�l��!d��]��T�=`�t>���O��Y�*1x���S�If�ȍ:�lI1r���9�9t�,��g�@D��){���=v6�d�y�{�D���Ǹ���x����>�憂*�ِ&�.	 Ǩ�	��N���ڍkUL5�m��c^��l-���"�������DPž�<`g�/������Xt�����8`��u�s���U���~y`�h2��+�c�㆙BuK��Y����ar��ġ�RVn�hv���Y��boW�&B�â���\h�_�����F�>�Q6C��"]�>����qH�NF��"A�ޝ8؃�ɶ�Mm�_����5�a:9)�^�J�m�6�{6���e�ҍ�v�i���5M�g�pd��t.Sy�*Q�2x����Ƥd�
G�};Ha�DO�Y��,��4v��T���ǝǹ�HD���eB]U#R�Ov�-e=�X�C���Q|>R��ڏ�D'����A� ��*�1 ��S�Z])-{P"BJjaZ�_��7���|r��A���.Y�X,��Z q�~sN0���\��}S;H�}��p4����C��	y��h�U��U�g;��nWX<�����2\{��4̙/ˎK�|�(����N�v0�� -  i�۰<N�}���#ش2KZ�;pQw�H���. ����l�cF��r��[{!����y��_̆�Ǟ����)���
4��t��h����x��N8�\������8R��z�(̪E!��I?��;�S�_�tn��_��l�����%:�Ɓ�k�X�>�A�a�H,�G$����D���.v�@��&Q�֭�������j_�9�1�D�%P��kvu����K�ӡ J-��, �p��m��&�ߚ#O�a��
	�`��!���go�O\�}�K��i���X஺.��$��=��$s�E�^�6� ��O
���n?tC��sh��N�t��Z��U}����%�(6�f��]�����G�Ƕ�H3�F�yWcg#�f��Ė�
�.��~���<��:�bj��Y���z�F����<K�'LK:*���惲;��qZ:�>r��\|��-J�]�0*�;7��T���L��ò�빢�pK�;<Ě������L���KG._$;�K����Pp?��k�������]?��eA<6tl���~�=C�< _^���2�~U@]�b���9���޻B��5?u����  `���K���5f6����5��MQW[�u�b����Va�}u�W�adT�C��|���H����hc�wX��N�7��H�#�{�	�R0@o�G�A@ޓH�rvz�����]4s����m�*�3A�L�}��g������}g�v�|l8��8K/������7��~8��,�4i<��Ł��.r�#���B��0^~�)H�)�˹��!	�3��|�l=�9u�C ��3���7R���:�\o�����t��]~YwH�&�����N���+^��o���N�:/��U�Z�R����&����>Ho�Ϲ��-V����*<�$Ќ	�H��w�ȍ7%�;�W��ro���^�;h�������εҦr;�PG$�#E!�|v!s���K	����?ݒ�k@*�53����*N@dy6�*�V��iK�!�L���G�L�r�s�ʢ��0���U���&�*b������r$S0�2ޑ�Gwa�CG�C)Gw����p�z��u^��]Le�[ր[��Vy�\Ck$[��E�ّ��� ���T�I��q�5�n6
�|�tWP���n7iA�hɴ$��l+�F���<��hm�n�"�DX�Z$�8�7阄6���M2�S�2*�q%�"9ؖYr	@ ��&_����;���9n�)��Z_�	3R��.�u>�D����v�낖��Ot���h�����^$�[z9�.�8����6��R�KU,[��3>.&�%��������!�J @:�!��8��_��*Rc~'��Z_'��}�)�Ρ��ϳ���T�0`)	j�ŵ��^��"�j��u`��g�=g�(��lYGpMR���*u��#P-�����Q\����.�8k�/����#��y-w�Ќ�dwL�8�h��u��?��1~�z1�Q�Bɚ��Mj��uR����	'D�  FA�ä����I��v4쫫�M����5�ju eB������L��0�웬h���ڧ\U�����s��D�$��$;!δ|5�����B�Ǫ1F�R��'2iJ5w�=?2Q@��������BD*n�8O4�'�r	}F���ыtm��]��V����&Z�X!�5�P���ZƆ��8s�3C��G��ztJ2��[��a�H�R�����IG���n��O��*Y=�ʟΖ�cL���=���ug��N�MU�D�J@`-���%���m�����)��	n���/X�IM�2۫������L�L��˱}����ȍK�⁏8�ۇm

��7��[�`����L����ʺ�N�y�}��;,0��k���)�IRH�s`¯�N�-�x&�"����rﮡI��`���>�*�*�N�fճQ�Z����?Q�?�6���x�'�[|�ɴBxd��Q�Qy-�7m�����������ye��? �σz`	RJ�.���I���{R�3�1@�*˛��5>zI��S�@_Lp)�q�Pf+�^�Bͭ2zr��W�G'd��<��G�~ܶ��Uɍ����	狨 |M�����pX/s��{,�����3~�JvE}�%��u��$B��~� qe�FG'���t��S��\:'�2�/g���Ѩh�;��������x�Q�)��T��E*��:Q�is0��&��e�����p8�̤yo{A<Țږ�pA=��;/n+KJ����KV`O/(�⓼pl����N��j���l�hϵn.mǥ����Y�˼���O�B� ��hց�r�,%	�kug�+2����ZvE�[�>��D����EЁ�4F�k�e��� \����w�k%�44l�� ��O��0T�H��Ŭ���:G���o%��٨@?	�-�dfZo���d�6�!�.v������-z�1��u�a4��ψ���	b��|۹-2���m��yTL��)�p|�0,���\�kEU��\��l
#`
�(��6-)	ӊ;��o�U�K-P (<G���