XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bޥ��,��Q����b$H	�Uv*�K�8<$s4�v���fK0�UK����������+y� 9��W� n�aq�cE��� P"5$@��t��p�NΧH�Ĉ=t��_Pgb���(��>Anq�~���I>����\�p�4@�&�R�I��������P�rlk)џ*�b�&�[�-���ْF�B!6��c�Y������u�ş�� ��lĦ����z�Q�Us�g�w�Ƨ,�d�ds����~.��n�w-hUZ����2Lph애������Gf��K탮�?��^�cB�����DmJa�ܭ������u��w�=e��U�/���k�:���c��.ۘ�r������sEs����w��	�Q�BQ6R?���q����A���`5�h6O;������-�GB?�cU�%h�O����e��Я��@{�f�q��(ᇵ�?'���6��Bއ�~ө؁.Y���~���خ~�<��>�l�B��9��O�CܠfT]X���L��N<ù9��	�{i�He�D�H���f�v��-�>������Ǎ|���X�LH��$����,��m��2h�
D^0�X��yÈ�dM2E)�E�^
�R���P���{D�t��BiC1��=��=�Y�(�A�Z����(t��;q�}U�;���M���5��̃(�X�vq�ɼ�����a�7_��z�	����t��,|0�-��2~c�a�����)`�X�$�_�rD%ڠ��&�Ě����3�����YXlxVHYEB     5fd     210�����D�A����0���VL$�7`��~8vvR�M��@=�SX�r��$
mI7�Wv�ۜ�Z����"ǐtU�E�P~��#��Հ�:�dL���5F�P���_������sQ	���)���R�z�� MEeQ`�@��We�~���$��f'2+����~��L'�d&���*����w�UF;v��B�|��y?دJܘ_P�ʼ�Q�/�KfJH����4yr����F}�Ahp Uz��O��"�?�"s*��4_Z@d�RyS�B�B�A���t��t���%�ec<:WV�϶����oP4M�rV�q�{e9����ʏAjZft!g�م ���Mq�3#�lAS�6��A�l>o�|B{f�HH���cPIq��VKg[�}��-_�tT[�����]�-�i�v˭�4	������sa�*%�9����r[������J2�P������A_���ϚOz@��$�2F����$j_�b���lS����G`�M���f�T�	G��