XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����U`� w:��,���p׭�<����H��n�0�����ROu��.���F��6���j%?�7��OA��
֔�9��J쾗�%e�<v�?�Zke�L�����gI�˿�����:�0���!��/����8�LZ_�(�h�]���ڷr	�F�/�>LB���%���N�C�)~�΀���E�-�X!�L<���`�*j��j��:���- w���W����ɅL��d��oĚ���/��$�+] "+a�/�]������Y�7��N_�Ƣ�TW���ُ����?:�;ǽ��h�q�b7A�[O�|U�l8�ݕ\E�1+V5B��h+j�x��5LN�.�	3�M�,��I�������x)s�1����C`�H޼<�p,@�OL'>����b����̚�|w�O<&[GS^bx�E�1t>�I�qKL�$ ��\���_���V�>3��$�x�A� $J�%꼵l,��g�K���"ya��e�̔�����%�M��œ	������X#d�j&�bzC9(��ro�l� �P���7��R�\��Hw�خT柊L�^�� ��<�2�,�T�/�AJK�n��d
j�������B$'�x�4Ga�ӯ�[�x�0��DN;��XX�{
[���>�7�Xӵk��JF_�O�
�a~�����A��P�Cr���tC��~�'���u�����*N��H�����1�A"bم�N��'P�-����7�ޘk�� �C�[-u����MwXlxVHYEB    5be1    12e0l_�&���?a�P�GA(4A����7��j�D1����ag~�>e������w�ܐ㴼0�toS�O-��+W ����j*�.7;���|g���d�-()L9�b��dW�<-cM���o[��:.�gC�Xo��
^��H!*C�|Lw�Q9v,*��10�g��5���U������ 
�ⷡ�:]�zlPnpHw�f�;Zh��^���F�����A-ц}�F�	�Ĥ���Q���2�C�z�����>"�Z�^��^O*��}�=4��*R��dݻEK濌���]��G1�gr0��ѣ7Q�m����[Q!�K\NE�c;K��2a�ћf�i��r=�Y	�7���Ɇy���t��
�7�I��۹�z�qr��釘fTؿ�)�@��~Z*L�n�`z  ^�C ��V�щ�$�ʉEx���F�n&[C�p��4�j��'�E��Hmf�Zܺ5<W�!��@f[�vO~g�2���2��2��]�����o�d#{�n�`�x)@!�M�(�z���N�|�k �Kz���J�o�&��ԭ�Qł�8����m;���깜��b~K�}NA�/�Z�tZ�x���k{��x܇���fv|8\���?5�O�e�"6I:��6�ъŨ�w ��څ�!=R�����t.�</G�lBFsM�5ӻ"�fr_T����LI2z���
5}b<�iZ�G�Ky\��O��.��i7��a��$����/�����L5 �-��>64f[�?�SD�]4`ݤ<cO}��u���=
�`��TԸȁ+� q��0�d�m�3ɒgc�u�Ӛ�GEv�� *䷔�'�~0���Wq=3e�~������lJ�ՃS�c�+U9Zɮ�e!Q't	�Z�;& ���[��[\����V�J�2���I�> ���:�SL&�P|�~�<��-y��$�^�W�8:E��?�݊L���Hh�**\n�a�E��O���ɤ� --����5�6��j"(|�e�B]��������R�y.U~ ��rt`X8�f��F�p�M�M�|�d2;���� _�3Ƴ�y��IV��D�ƀL&I�����c�����p���Y���;�����Hū�|b*yS�����=C��!�&a�?�nծ[��1��_�:��l��c^*�8͗�F�zu�*CBH@�=�Y� �P�-�m�x9KG/�6�����ڍ�3�A�t�}H�=�a���ۮee�P�5�'��)���`����;)t�p���sl�Z^�J�!]�ɱ^Ȧ>>j]D�q��ײ@��R!�uڀCW���ø��Kq���8Y��Ԩ���H�}b9��y
�����-!-���b���R``8�ܯK����7��4D ����"�]X��2�)�0��>�=��[F����c@��đ꺜B��L��xF�$��q��bl|]������~�	�X��*����|hp�$��ųW���@J^�_ysHj�yOz��U�>lV�S$��v��}��*�(ܑJ7:x5��X_tUcS�{솿��Xn"���^d����$�������_M�����]!�%��~{�;��֜8���S�a�}����~��vHG��7\����mta�%o���5���x�]y��ܶ��{4l-��܅Ƽ_��G:"Z1R8����,u=�6����,T=J�'�]�&0c�Zi8������1�;h<����W�'�!���4K:����ܺ@�|aB�N�!�V��c�ۍYݎl��g�W?#_���5؆~�R����$�O �l�Gɵ��Yr:��oYQ�`��y�� ;& �+�ط��f����p�h�wD�֋��u���/���������@ls��d7(ns�XU��]���8�a�!�@�F�
v�u0�7J�Ɔ��w�	�e1Ne�C"��rE
sE�����5Ȍ��wS˫�H]�b�LZ���o�a�n>��mt�.��'ŢPx�x»ͮ&w��%�A���L^;��Ͽ�R\�`^�t%nm�ݠl�㖼(Ѩ��5����E�;�-B�I�}���3ow�n�����F���a�UKE����FNC���� ڙH���)�Y%��'��,m1�݇wyo	���V4�"'8���K-��$�8�Sk^5� �D���(�>���I�L���JkB�=7TW��k�� �^�)rr�8P:�p۝�	�ȋ��{B�4X���5�>B��kö�a`�6uze����y��)���(��t仐�_��Wf9�LI�6v��|���R�r>�#�NVO�� ���<z@8�����Ub�����m�W�k�5O2��i�u������^Y�^��:v`�u�-���)���ǝj�q�\��7��&ĩ��9-{-t���%4����yǭ��4?��W�?��AS%��؇��Zr"�[�{E��6��E���Eq����� ��wqXpK*+̝��)�7����;qM�q)F[3��6���S�ˢ��^/lo�M(�Y�̛Mɛ��G�����*{�_��~q��h�Z���ϵG�>�`�ؾ��&��V~Y��t�^���֐0��M����4�Πa7���࿱��7KW�s��cЁ��c���`��<)��i��3��K�Y|:N�]Z�EF�[�Y��Z��=�^�G{ �H�/���Џ�tt����»r�ȓY�Yl���{��8�_1a��}���H������B>P�]*%,�:�'��y¼��蘙�b�qޣ�@�PG�F��p�͋��C���,"��lG��ΣG�$�iwF�.~��:�6?��m���z]I���xTnң���l���#4��Ҩa~O�hUI�?G�/Om3�9B�g����$�t���}���9c�MŁeS�SE����g������ae�_�/a��俻�Gܐ���n1(趘w_���tJ
y{�,��q�b @ɦ%ż7�F����."����P���Bܭ��Ug^�M�갥�6�v`�P��҆e�&������'��:~�ܽ����֩�!GA�����)4o����L��K`�h�']|ӱ�M�:h��y�p��+Z}�}>���IV�e���Ƃ�(X*�v��$*b�����n���䌽!�`b=�D��"�IZ+Մ�������p���
��!8�2??d� K�Ɉy@7��\����9B&���a#C��{�@����~�<2��M^�]���e�U�=������#J�yq����!�j%$���ZZ����߳��UC��1=�eS(Ϭ.*b��lJp�R�a=�g�CB��2Jq������H�xW�ego�ΖP�0���#-�SS���N���~���e���>~��O��SxL�n,Q}��߫"M i9�|�N���dQ)��E��Usm\k$<%����ǵ�(�;�0�����#v����$G�S��|�N��l�sY&�,� �f5՛��\��6I�L2�~7�o�|���F.'+��~mUPh�Ǘ�-�E�o��R��#]�>8�� '<Ekح�}4,1B�!<H�Z^�-?C��z�bw���WA$l�"�����~��t�R:�Q���,>E�ʥ��ڑ�s�g�ޝ��m���>�0��E@�s�M��)U�q�����hMj�xD8�3�z�7����z���g�4s��D��汻\=7�]�Y_��as�=ص��n 5[]���,�a���7E[���C0���/� 6-�1��,���!|/�e�~խ��D����� �{,8 ����+mOK���3-����98��0��]Jv�G8�w���.��P蹛&}�������ܵ=P�����ԹU�iN����2��6����Tl�F��J�H�EU�G����D����>޼�,^�}b�eT�л��ܩ���9���$���ܡ���j�������씧�{K�]'�f�=.6�� ��#�"t�"�D/"UF���hŞ���*�%�싰4�|c��K ��L���fzp���!4H-e�W{�ZZ��k��u��E5%���F�����dR:�����Xy�r=׃�c-��[ӿ����{V�)T!ڠ�)�����[�����{�0t� y���b��x_ֶ/Ћys�E�C-ĉ��V.�j�)�@���Q�g�_�O�%(SH�
M��%�Q�� �Cu��h������ڽ8
�ۮ�5�K|��R��#��N ��Q>v���$2��&����|2��Sd"9T�ǃ�q�lVA^�L_]_T� >*=|�q�>��$��̄�4���6@"i��b/Vu���}�,_�nHU �����S����=��Д�X���U�R[W�/��?��8��H[,<,_~|�%��B��~�Fٖ4v|��u��+azE���1�S�IP���7f�A��M��j^=���>��=����[��|u������ԥ4dA-W�U��#BQ�>)�E���]/�H@�]�t��!��j���]#O������q8�.up�I��0yE��jw�b��Z��?T�
���$�E�%�_���P����8���f�b��^T���MR^#��t-��G�����b7��p&�Ԟ��`K���K\��0���I3M���P�kX�Ej��Սv?��v��gv���`��������Pm�s���3���V�4�y:&�HZ�����K�&�l����x�_^���s\-�{nw7,������YAI��ϝhT