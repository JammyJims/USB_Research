XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Yr- [�+4�3�@3�.QƆdC|��؏��nKC5�e
�F��<A�r�r=S��� "�`M)�%8��9��Jo�vĸ�U�;�0�8�F)xj��[��*�pT�����
R>آ�-Wj�$�.�X�#�楬G����;&S^��>��S�y�FTH}*����ȡ�R坼��MXYR�����f�3���i��E.}�a�P�A���!,D�h g��&8�sTGU�pHٝ�O	�r��;�qʦ�W�z��`o}��P��6;Ǻ��*Й�U��y��Z�tl,L-h%@�2,׾q��qg��:}S/҈0�W�A�+�Ds¿����ɶ,�	[��ai�iV#�H���gU
�ub$d�J�/�59-���]�][~nN%�,��2ұj�u(����S���� �o��&����鑭�}����ɔ�ٷ�J_ٝ�	��>,�����:¿��\:o�y�u,9�u��r!g�L�X̍Ce��5T-��A���R��~�CɨW��������=Rc��]��x�� �{�^��aG�]�Ż�! x�>ls�����%=}�7�C�572��*�c= ����$9�xO�����y���ur�t��'�۞�a�1�>r���`ȠZ�C�n���)��$r@�q��e��[�c�=�8o&�&V+*�]�vc��3).�D]agz�YP)��n����W�e<胵�J�R��V����:�13x���6D/"��迎��PZ�Z��mE�5Q�G���	{XlxVHYEB    40df    1270#��'�O�.�]r�8�xf��o����3W������^b��a�RMѺ� :�r�zx�p뒡��Q㓪Q�;�Ȕ���j�R6�_ɢ��>\@�Z* F4�o>p/����A�)T,���1+��d��Ƃ����ٺkYh�"���q<Q��H�o�r���{60y������Il���ʪ��|Puq��J��Y��N��� ެ�L,Qi֚y}ĝ��Jm��)V�C�X��Yh9��� ��"�u���8�Y����Ko���o7$/"um��&@�;��*�@Nh�I-	v�=�����v
���g^x��6q��[�,C"T�%8d )!�Ci���t.�� �s.�������tֻ@0�<���)~����0��ђJ�Vx�]W M|�7��Dҟ��j���e�	pk�
`�����v.���$��(��C��G$f1)7O���i:>�UG~��P�� �ͺ`�?�%�����c{���Q��[�/H5���X�$3�'b\1%T�Xд61�rv0e�c�mO�tR��!,�7j�/����Ԇ� x�*Ms�,�)�ԡG���\�P�����\�>��/X�X�d�ʻ�+1F��}��s����4��)����0�B�Ȁ�ј[���KD��<��6�E�d�*�j��z�5�;�E��v W�� �ʏ�0�@Y��ʰ/c��%�0ٕ~&�8�u3�v������Gn3��yJ�p���r����]��8�n�����>�v`*=ŗ�YQ�˦;�b��ق�=��nʮd��$7e������7*sE����c��Ǔ���
��|��ϷCufM�:�:�T�G���R\�s�x�)�ь�G�L������HV�Uu���O�^V�c����\��3�46/Q�����釘�V�F�d��'���R`����|�k<�mq[����i�bE�@��:h+�U�IC `�6e�B��Ͻ��'�#%m�6����G���� ��Ĝ:կ����( &���8-���)5i4��t�)kxjق;��`,G4�ɢ��S�O�efţ!�L^
�0-hRU;�7�|E�&���T���AK��� }[�3��n�|��c�ːvꉀy�x�s`����sL
�W)�	�k�?��*�fPX3{�e#B�)tUj�9�G��d`���������߂l)��S��B��yGs��:����4��7>`����DF�n`�h�,Nn>��!/y����C�މ
�M?���v>S��a�1��M��Ŷ̢ʡt��U�5��	�U)�쓈���V�8��Hնˎ����v?��U���x�P_ʫw= �u�T�R
��e</�[ƥV��u������������p��!6E�l�W
�j$��,;\��L�P�e�ӎ8V�� �R꡸�L�ETd� �F�L5֓6!b9�A*���n���� "�ą�{�5�[B߿kغ-���),.�Ͽ,;}����1E�Mz	0�ݒ��ؠџ��/~������)MD��:��zP��ӏ*��3� t�Y��&r�"���5\4���w����=U�H��y��5~,Q`{�*�V������@~�I��J�d29�{����̎O��>����ۗ)��z�����_�(���ĊEyڕ�����?�kٺ�b�G��Փ�k��ZCX��5w(�6��]z)Kd1�������!��0�-�3xC��e���.p߻��w��#���p{�vM|�	�]ݬDD�pH�N���'p�=� �#��Ԥ7�.O��,9�~��<K6��Ƣ9��Ħ;"���Z�D\��s{"���%i}H���M�[�&.q^�UРk�a~�-2<�@vH�eT��>����s[w������N�H�?��/)��&��{|�2�ZG���'a���9�x�Egeg�n9k'0�5R�[��+cs,���2���"r��CS*�L1r�@vLBJ��lf��k�{3�3���A&R�9���4-!�]����t"�	}�oA���P�A8���)�#�c�o�:{���Y�J@(���#mn^�-��������ȵ�C�GB�k5P��6Yb�߳د�O�Qg�$�x�rg'���G*ʽ���dlV�~Fe�vW>�����@r�N�f� �QȆ�x�KB�<GC9����c� R<ئ��u,�H�U�܀�c�g�)�i �s���$	~��b�V«��id#�� ��uz3#s����H�lw�1���q	rܺs9��g/6�v0pV��I9]�=X;(-4ak�;3M(P�+��t~*����v�ZN�|����5�_[ʋ��E8��YҎ5�ȝ�C�$��܈dI���L}a3G��&ٽw	%`V��MB)���c���;�в�'�T3�%�&�'3oF?�v�bV��e�5�/";y�$��*L�Gw�1&O�L��p�)b�\v:�(�Ѩ�h�"6�%�=c}�R3��ި��R���FU��/���I�4��~3Y��Vq��,�J�k����@hk�-MlK��(B5:o�� Ұt����B�T�9����C��(��x>��F�c_�m��T��s�j�t��#j�D�4t
�TG�8,�Ü��+���D��UZ2��䧙8�uh��a���RH��1�7"���8����>�C�#$���ʫ��H�d��Kx�����v�W�ů��;1ɟ�b�����_?U3� �9���E/�����ǽ�uk�x���g�9�}�^
�YAp�A��BxDd`�$�{�⬬��������\��O�:��Yv:X��'N��,]�����<0tq5yeeQ��Y�0Z^Q�t���+x0�kƔ����Qu�9Gr��RK <�LO*m��Xhҿ��w���L����ε�F#���FtDNE\JX�~ҭjw�[��|��c�E�֤#�\��^��y�=��]c����9�l��re��4%���F5�"�dĝ-q���D@�KM�:�׌���m9q�����e����u�&�9�����h�}m_�`�����?T7m$WU;u+3 �/�a5���������@U����Ct��K6��ɇĥ?{��,"D��>N�	Y�I���v浹F߃>��ѵ�h>���4n߬��쨼J]<�4C!��kR�9�|ejJU�_�����x�x@H�����d����W��8q��Y�嶧�>Z8�;.^�_��[�oͧ$�g,}��Qg�Vy�$��)جbOVË��z�����z��uS�c�B���=��N�B�޻��]||�U�b���,��o?��z����CN���[b��j�D�.������p�]�lY�O����^�>�s�v~zL
ߦ	u������cwQ��r��@�֯�����4w���i���Z�撱�>��~Yi��e�� )�f�oC�z&�K#T�:�O�O����%q"-��N���$\�@$n}c0��4Ť�R��=\�t�)�i ՟`�p���=��&Pto�-G�
,�A�B���á����G�������S�%����ƞ���o� ��k�Ȯ#�mo��R�#�ᾅO���̥ԗ�r�t�$z��0n_����j@<��������w�W&�᲍�Qg��c��d�J)�a�y\�#�m{'���c�D�ؔPha|�[O��f����xm���CG�e��nr;��*Y�[Qdj�>"���j����I���e#q�+DSաi>�b(:cEm�R.�a#��l�21�{N�Q��4���4_�m<��&�Uh��*ߜ���k�oG���3��EvQ��	Id��x9�6��ТV*���/=a�n����Lh5���ۚ��TL��>N&��wSN>����'���ojU�f�-4&����RN����t�;eٰ�����aDO�=!FӴ�T�q��*�5*Rv[Z�T~3ܼ5ϵRP�ħjQޜ�Ě�tŕ�X6|�]��^�����gј������x�1��o;� S2
��B	�!�Bso�L�n���0��x��y��8q�9��]�~�e�b���t$���L�q�P9���1E嚗-{���d���[�hp�~,�vm���c�D|�F��j�J�r�>�3�Q_���@�dV��t�N��#������ |�.N|�� ��S��줮N�����y\="��S�.�{�_��W�/�D}M�O�O�(��+�]�Ռkk��:j��CV��L��J�*�d؋I�Y�i �@��V^7��db�]R	�������`�Ӹ�2_1Z�8&���i������jgq�az��	�k����٧�����'���Yq�%U�l�w��?�/�h�������.����|$Df��^�[tG�[�������e��,x��@��WO�-�m�.D�S�{Bn�έ���ie����� w�n�}�C��.i�@k�zC���D����~E	@9�[ba�_P���~�oz^Lv����������Qtz��U�I����K���Y�V�ɨ4��m�8��>{���78U��+(���V��[�D~��� Q��@�c��u�(��ֿ�������!=D���H���+F�@z��q$��^�c}ڔ���2��o�м|W9��t�X����v@�T��'�Ӎ2