XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~!)p]㓶V��8�v~/۟i�T���PsH��_�m<Vz~!N>s/8P=�$	Ƙ[�}P�Ⱦ�E`1������ђ	��T��L_g݉���7���X��ry�v\C�HVa^AJ��F�r/��MlO�4ʠ�4��tUgܫ�	�^^Lsgi�$~�͚��:��!n;Pa�*W﯎t+�w��qr�:3&4���/��<A8�ڬ�2�}��nE�(�#񢌶�� I���KX�M=��:h�X�w��@N5�|�P�1	�=T"
����i�U���O�%��t��t<_��/[��m��lm��M]+t �Ҥ��|������ٌ�bx]֜7-W��N�YD��}�{��������ݿ���P!�O�Aa{ۀ|�H:����F����Ẁfވ�譄c��F�\��u��X",��RGh�9���mګR�B4D�,[R|�K��X��K�Ѭ&h�,m ������C���ߡq�E
���|�;m��V[ h;�z='��礰5~9�;�����hB�:%m4�6x� ����l1�/�2��mc3O��������Y����T�����m�N�J�S%���k�l�>�s5�-�B0e@�o��O�)XB����i�+�Ӄ�[?��+&�Ѷ��F;�V�H��������q����:��G:G�ĸ�P廦_P��`�pʯS�.��{D��g惆V`�}�i' $�7�6(��ڴ4���GWi�Ã�x�H��t�=Q-5���F��Lݡ��>�%��^XlxVHYEB    654a    1390��N;�
h�tg��7k��_�$;x
�-�w��;��p���&�F�h1Br�ĔpRX8���!|�u�%߱�`{��1�R/Jw��)rꃥ3�͚�&�� Y��ɼ9�dߗ���:Gf���J�a\���ef�����ȣ������S�}������l��s�\��'��h�M����l�ҡGq�9�_^(�qZ��YԀ�M���3)v,���L�꘮ȩ�A��'&��_v���
�d-e�e�(�G ĭ��x:��n��R��h`3k�1CM�����;����<D��^#ȉ�f�"�(��c'|}�b�z�Wf����=��!�>E'���� &�W���~-���'���E ��.t��D����F�b��ȳ7F~�	�q%�5 �����n�N?z�_J�!�7
P��ۢ��}"����F���H9�&�,������IPv�%�'�W�]Rl�nu*�~��&	LJAta8�^ڌ��x�2���O�<*����<�1t�|�3��B� ��3�Ǩ�8iZJ��.,s���*J�����gm��a���9/�3��TK��\|���'�9ѨI֞V
b���x�Ƙ;��\D���D
�GÉ=@R#��+灘ښ�C��/lXo=	�)��Կ�b�UqxG�({�e��]����}����]��[�|^��o������B�`���n�zI3�^�w���8����s��St���͊��b:�E��#�rF�I-M{h�,Mօw}Q�I��J|U�_ظ�ƴ$v�ޝ�����P�����J��ܸj�7x؞9��\n#7��/���:�H4��_��s���A��w��0��Y��?�Q�I-����� 2gkl� X?za�<$ ��o���}��i���D��P&������h�怣{&�_;f2N[,T��K3-��j�W`M�z������qbX:@G��E+�����)|d1����k�Bu(���u}pȖ����Q{	jSOPo�I�#,������~O�Br��u4 ?�*���7�`�6��$�G$$����K����F�|�Ǥq��C�.0��ն�F�I��>��Ma�t����N��e���+�C�'���G�Yn��$�z��ym���D^�>��ت�B��H
{�;� ���>��A��".S��z�IG�Ɏj���G�}�<�4�P,�V٫x�W��/����ƟzgVѳ����k���2��k�/��{��e��Zq�����_�����[�%�>>�n���e��hXS�s�B��.&5��*����&]�u���	3�NVԮ]x�/�`�H6f��D�g� }$1���7��N)p�c h� (5B���+�j%�s��u-����_^ܬ����g��F�>�:�z���g��3�D��yF�0]�5���f�h���0N���̄��r���� Ź5��
�t+u��=m������u�l��R8�w��M���{#�F�]��̩�xp����S����W'F�S�Ţ#j���X&ms��a���asK.S,�?�ݏZ����K(]~2^JW��V$G�m�t�*}T}悎�r��bTU�T(h(B���;آ/���B�aуO.Jl�}:�B��z1j��[Vp�r��q��_���Ƣ�M����?�B���� 2����>Ȝ�<27v��B[�^�\d��u���o�{��A������v��B�҂�`n�zW)�(�a�c��{�����R��.������̎�Y���
d���oeE�k�C�
�懾�==��! �tX��}&��j�=��nM/�Wl/$���E֑(BE��J�~OK��"i#u�R�*Gk��?��H�X�Q�D�AHǍ�%��/C�꧿�r�~k�y�&l*��5�F��"7By�|0��wc)���*�J]af�OX>�ڝ�k���tuDq�d�ʖ�-�Uɭ��ݭEt";��Ś���6��9~'�F.<��L�m%�`��k�F*_�_=�K�8苩�4��:��c)fa:��M��m�������D��L�����O&ck�)��%��9e˷֐�$g���@���i����|��T�Tk6�E���D�IJ���sD�/h�4�~����#Gm�5ZM�qXT�c���>B���;g)���b�����5�k��)��������<�L�ZV�^��d��C�G���*D��H�wq��P�)R���!s���W�Ҩ�e�F�9*Bɿx���n0������f��
�I�3-J�2T�Mo|��L�	�� ���xZ*���+�jm6�T'ZUX̤�,׆������)�.��Ux��s,W{��2�T��JK��N�_�н�p2���q�@��!z�ʚ'_�Z�7J��L��� W��ܜ�n�Am�>aP�����q\��7QZJ�w�tP0Q~e�뙣|�5
m�p��=JQ ���خ��ª�#H��}$e6ٚ�/���`@��E�"���M��P�d�u� RZ�;��Yِ�t*dJ��N%�Y������E�ʺ>�c�+��4�Zt��?4��V�n����ޖd ��1���f'\[ǡP�Q����͈ ֖��P��iP��QI/W��H�/D~/�H�~�.T�YˡjG���령�� 0�,�$\���&�c�ʏa^%l&����}@mu��Y��pF�=Q�����_�����zvc���@
��l���؎�pt��b�j[�V_+�-&�ڪ}��R�i��6?�3�M-�L���5�ه'9��}7��b[���Ӫ�B��,1`,��*���'��jq�ң�H5����#�4���,�xfU��B� �Q:)X���O��rɵ�oN!�DM� ���h�̂�	�||��Y��؜�7��Q�WgRj�a.�N\����)���gA���Cr��*/e�	A���UD&4ږR���#c���!�fQÃ�pe�M}�xzV�:%JH�&������世���{�z���d�RR V�	w��_�&���vQ�8���a�HM ����/�N��|���P��?��Z��iXkW���jz�퉻nu�<~�XEx,ѥ�8.�(a���\��U�.��D�!Z�&NP��i4�!�Q��F8�_�K̷�D֑�g�H��hv<�l������uz���W�ͼc��nFv�@��.eg���]��]�ba��7���gYk��o�)w�z|q���	��}�O=�r�۞��/����h���!64k���4��0�$h��.�5����<��I�U�ٰ�/H��H�YL���/?�q @#�;�]�T|{�鋯9,5�5g�v��A�����9��0�yl��	�QЋ��HYz�&��m�c���|�|�1j��cAZk���J�o���Qg] �ìߐμ_Ţw�v;�%í:u�'V����TMn��K���*��Ѧ#]�'�G"?P�Ֆ޾�� ��c4[�+$�>9C�1�ר'�n5��h�����?9�h9ty�X=g]�17"$}��*��E9�Nk�P���l�'�9�K�Йվ7���1�5����/�\rA�@@��e���]��( I�e��CaHd Awq�M�|U)����ܵ�R�eM��\a��h:68x2�tM�SJ�p���zp���	�'�n�@w$:���0���B�\��U���޻��"���)�p/�3�1�#7����H�a�Ѳ%�co�<��t���@��E/2`�*͸ϡé��P4��㤈J���|`[ִ�}1DU%܈��\�f�G�˦�CI�`w9�]w�>�_�W�a0/��ګP��)�?4�Z�Z�p\���:���w�_AI�p��x��ߠN#���U�;�h�����ָ�q @d̉���߇j���0�Dϧ8�R(9y@��}�K�R
��U�$g���nxR4[��O�P5�r�����9�	L�����w.�<����2/:̱ 6:��%�Am�E��^&��i��4�4���:O��'�}J1��8Y�KР���)��fݹ�aY�a::����$�3����p=g�H=^�,<�h&�$Q�#d�~���_�}JJ>9D���˾Z��ܥ��Z���7J�#�C�V�VT��:�	-��ݻ�Є��{�B�N7�Ӊ��p�`�t{���t���]���~��=�z��O�Rf/�˧����~J@� ^����1&P�ޡ��u$���;�+�HmZ��XI+��Zf��R�ch	���ƻYN^�BtTcs�:R�.!p��s���]��#o?]�f%��տZ�j���T	p�⒨R5_-�|a���4g:�ӫ$͎�i�� ֬�]���\ԋ4�U
�Zk
�5�o�)'-�|%�ev@����}K��3V����ʈ��'I4�P>; �kBrR!�6^fT��q���J���K� ZC����9�n�A����ē1mHL��GP�u|B�=EpLYm[Nr ��R��(��Z'�?	B'��5#p�Ӣ������*7)o����D�1o�ִ���@˹^�����|�]�t�Y���d��n��dEd�Հ�K�ǩ.�u�����f�o5��bt��.DpQ���F�nᶞn7��XY��Mx�X������[/.�<Ν/�6u�p�S���!6�ƤA��IG��G���=��H�O@����;�5d�����:Ů��k��Eΰg񢱚w�ͺMEit����;��|g��: ���C�� �F.a���O�e8���je����gp��]��$O%-�.��BŌ���%QA����6*�ۛ~#��4@�-m�e)���Q�S`��֏L����%��qBClo����2����Rt��[m�33�tMp��&n�@��R���QW�\U�5v1�
�Cu�Y`#s����}sUs����]���/�O��� D.L���v5����qTՀ�����c��#ڪfY��c�'�p���(�f��9k�(z��!ΏoD����&� �xJ���