XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�^?T��5[�@}�\�`�F�}�u�/�_���9w;S�w��HPc��y��ʗ~Y�/��s�}/��ʳn��(�v�R�[W�.���!�߁��6>N��λ�ۅVǚ�� �w;��z�@��l%8��b������ʽ�כ�	� �D�;��x5��bвR���᜔�/��%���*����|S�cTX��cx�ɰѳ������o���YO[k	_l��H���Φ�������~E���H��-f���.�pz���x��[����hr�
�=60I���ѧkS��w��t�C��|ϰ�|�H�ČtU�OE'�"��S�+�]��F�7ʶj�%�ueΏ��8�l�c
N*�f?�\�k��bU�Gze��/��\e^�m 9u��?ƣ��\BhȨ�d 
% [6���� 7��Ԉo~��>����PP�Ŀޓ:�cG�͠>D���Ud9UK�^�(O�fH�g�����F��:�k��\sc����JzHîI��f��y�m ���4������\m&��\���3�� g��t<6��C��~�p�Ku��6J�c���Rl�%J/����¶�����er�QіGb��q��&�Mq�^�3��MjU߀�u�Yt:�dUA���zN�_)
����U��@V�F5���V9jb�=ݘ�_���7[G?j<)�TS>������c��;ΩȺ��� P�?	h}�c����:x�
[ZiXE����C�j��ʘZo��P[*6���XlxVHYEB    10fd     700����Fz�j�Ѳ�T���G�r븼N
zM�oi"L�f���/���u���_�������6�� ���FE'U�	����87�k�煯���h��PL�W�_��w�JV�Hh��:f���!�X3^�I�-�����EB)ST54�<�KX]�Q��lg~�Ɋ���8Ǉ&�ZR~&��FU���Ȋ�ٳ�&�Z��/U�Q2(�������}�B�}s�X`^�M�4:5o�f�8
�7c}㏸�bVQV��rp��cn�G���rL�L׶��@M�f��1���%�j_v�,]Ћ�S��|�^Vr�(u���G��C�H*!�3��G�Z�[�2{���C�1=,Y���`i�rA"a�/�2��r�9{�nد1�{���XE�i��z'q	j��%�I�j�dd(��B=��-l%����S0��&����l�Ԛ��p����F���A���b��i+���;�ynVO3פ����4R5,A?�0IESqn�����4D��E}fo��\B�ʛ�i��=6�)�Wߝw��J"Qݿ����.ܩ�r��,:�=�xz��~&R��!}J��S��fV������tM�Z����j��@����b��Huh,˺�<N�_[�m�yj�+ͥ{�z̍<�SH�d,k���	Ȗ@�B�h�N��.�.��^+��;��E�٣b�7����]t�G�L=5�K��_�6�fz���$3��G�zg�gRuk&'�O��T$)�QЪӎ鳙r���n�w�:��w��P�KT�+��ǖR.< ���E="����E\vu�P8���?flE��^�r۬���e�n���`��Y�eQZ���c�2|b�܂�Dn�p�03J1j)�_}n������m߁Q���|<@�<`}v!�)B����]�0"_��6%*�Շ�}1��D0��j�L��f�Ss�[)�k�<�v=h�]���m_��vcL��m�4��ƻ!:'j{��2�ؐ-Ø2�7%b�+�k&#y1ɣ��d;�b�?ڞ>0���6-�t���V'����}�0N�5ؤA/���77j/]�#M;$} ��E�b4FY,q���iQ/@�c�\�^�%��rU-��+��pp���s�ҫp�q�����xD�mA����(D,����`J�Ydb��d��WoWZދ3�OK�$��Pf|�&�9Q��
�.�c�
��k�Lےi�D[;I����1��^-IS�4LKq@U�<��7��'�Ƥ���TѬ`ה��&��U�ΖY���V���uvגZ��S��N	��%Dn��y�(�{�Sl�`	@��:@��^f�(��Xyح��Qa]�K���T�cŬ����J,6����C\��Ld𓈃�	�~�((������h!8�F2S<�*��������3T����&�iK�>��TߪY�*j
�����H�(
4�lD���Xs2�y�ƅ�����nw�NM�<�i0i��(��D�����-�c�7��ȊwNu�45�9GG;2}�퟼�&E��դ�=�T��)�����%�d�\)m�x��k�4Yo�NaH���oL�{�����I�[X �R���JZ6ٳeX� 0֏+)o��|��z��Tn�v�u�l�O���,T����5%�B�{b��'#$�4���`���� p�nf��g��aE�=�r:%�ц��v@q�0d���tl#+��%�듈r����`�����~*X�xб�7>�JT5�c�
���e'.��`�B7���kҩ�}0d4�{���j��N