XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J�3O�C�Ǳ�]���F@�ՠ
��E���
����][�U��,�l�Th�ihUHŰ\���"$�e���R���˧���`�FFP��&�]�u��?�Z=@,z:q"�M�����°!����^G��`
�f�:�+��E���x���r�l^��vG.£'�[��ݦ��ǁ�?r�:ut��u|#j}W���Z��/���6�Y������Q�)8���פyX��`n�2݅� $&Q�':�nO��!���p�:��_�����9���`������S�l��ɾ�t�#T���ũ��\λ�oqRFIE����FV��:i1�+�߻˵P�+A�G��9+2��ĊR�Lu�o�� Gr�T!6t
_F�S�42>�y�� ����vK%�(�j��_v|�]�ߕb�S�r�p�6O^�0j��3Ɉ���w��ۓb���:�M��3%����
����?��"<��}�����:�n�)�^6��H�	YݲGx�&�.�-O����i���-'n�0*�3%���Z����nL����v�?�=����Y�[����p�6�;����b��Õ�$/�p�DU�Rƿ<z�q�Ɔ���/؄p���2L�Y�6z�l��S������g���� ��K������4^��<�j	�`=�-���qz�NIբô\ao˲�Eʹ����C�7
�q�˝�	N .><�I�������|�&�Ń���Rv)�x���5���l��� ������XlxVHYEB    fa00    31e0�q���p� Y�p�
���n�l�S_4T��"#0���t���[�|V?B���7�Р���uDe�w��C�(ۖ���e*�":�mc�e��UX�y)@l�<w5��y\r��*1Tw��jV:A��=s��H��;<"A��HF��Q�X9S=�f
�ٷ��	�Q��^��[R%�-�a�9&���`"d@ᴗNT�q����+�<��-�v|��(Vyw��4@��9�ΡyY):��@O��<�ɹ-鐆�)�=���0�+ �8l�Ʌ�׿�*A�8���	a,��|/�e��&WBA��"2���y�c�p���o`�Q�_t\m�x�(�䣸�M�4`B��;��	��^K���|�D��"�䑳/?����̴�N�A�oU���5țˋN��@-,���1��M+�~ǿ�ޛ�mw2�zN$��������`Q;��ìڠR��+���t)�`|ֱed�Xhw9�9m+���<���o L�Sa���p�Q�Ff1:���ዝ���T>ߒ�� ys��6-�̣;�cs��g�p�s�5�������5�>Q[�yJ?�	��h����+HL�#�\�t�Y�@��@��ʰ�ٟ���5��r<2�t��d��>��W�"�B�L�Y�|�0�h�0~��{�K!�{�tڊ���M����pqb�W &�+�lL:��2CM,Z�j=�;%:�X����dȐ$8N?�]ԉ�M4멬���QO��|���*sҢ�3�O���#!	k��u�8֥]�c9��\��J
��*��ʅy|Y�l�Ъ�S��WY?���Ĕ�����*x�]-��M%�����Gl˸�a��d����#��/�]��ye�*u�eN+|�C�uj���!s��!u*��ù���&�[����)Ry@��%٩��"��%X5���`i{s�>K�6;���:Gjp{ʼ|Tl�Vw���!	�B�=�g����p[T�%~!�uI���1s���ٷw���,�o��6+7��e�aR�)��x�Έ�.;1D���A��WI��Z~��F �?����5Sfe���c���t����{�\���'�vԤ
R� �'pnd�8!������[�Tc=�q�}�>ōh�g!f���q�}k����HY�Q{���<�Q��/��Y�����QX��1�S����+5o�k�Z��Ѕ�@ʨS<4�g����94�^FYy�`dп�9��$~�,a�<6$&�8L�M��ձa_}���e�Ͼ�:��
H}��kU�/��x8����Z,5{?Į�~�k��R��qMQ[�xj��g��9���m�r���ZӊM�ŶW�#b�Iu�O�P^EՊ�V�˖�T�d��DJ��R���L�"��[���������;����c����-�Q�b���r2D6I��H���"�M�	q�o�A�\�����5�n�9�$˩<�'��V[q���+4u�r(1��:�IV2�վ�MF�+s	 Qb�IC&`�\�!盯]O,�Y1&k��V(E1�`g�_r��.%-Y<o��g����u���>���W&I�����+NC��D#q��
@M��	�U?�LI�)���F�KŜ�� �1a͂)�C�sI��9�s1f� r��������TO.e������k^�^6#1�o
��3�����R��A@�䵫1�N��ď����ރɤ�"ô���G ��B/kS9�،H{���c���=)���L`:T�)��_�:=�
ɛ)��</��G12�ک�����T�2iq�&3���\dKf(�VL*�aq�IU�fa:�+y�n��i����sB5�`g��,�ˋ�*����a�N���/y"����� �a�5ֽ_C��BoE	h��$+/�*�y�`�?دU�tgFF��&��$ahT?�M���8���5s5�cJ�:���xlB����Sb�m F�?]e�9'I��'W������Y���{I2̽t�B�K�N1|�!c3�����`jH��T���8n��IX�=U�w��U\�ܑl$����rg.��0��S�b���k� =m��t@VZ(�i����SS�\��7���n �;4ױŴ�`��`лy,��> \�f{�
�����c.�R��Pe_N���S�j��G�j,�PC�������W�bN�v�:%*�����D�=���5�egqճ�(L�j|�0��(�籠�4�ǳT"4lr���i����!0x�zj�|���%Y�*��!Ƙc���.zզu�4d�M2B:�v�Q�H��ۈ�k4A]�y�h�{� ̡����w�v�A�U��QBn�D�D��I{z�w�.L�p���\"|2VZtB�`��������D319'�U����q�]� ��D��
Xk��xc[Ԧ1��$��j���yx����&���m��?��V!KӢv�#ٶX=?���Ne����h^re�;�G�)Y�`cV�G�l8d�f쩘iYv_k�7�ȧ-Ѝ�H-l�Ѽ��� ���?�/z���W��ËP��=3z�%9_���@|�Wv��A�y:�^K�,�-"W��������&�G���K���-M�EFp����A��Ø「���?�6�[���."��U(m���Ea=Ӊ��	mk8cV�l���_����:�q�gHǤ(GIBx�k7�i14-�7��!�����܈�v�f�.&�i<��>��2U�O8�V$6��E�fW�P\����n��aR��)�	��.BU8�<�N�M����H�]mf~�5R|h�4������P����:2!�s�����ˊ��E/���~<.FU�*q��һ=1��:`�bo�[f��5wkŖ�g�����L:m�n�N�Ύ&'_�%a�liS��\Ax�%�G=y���FqS��QַNЎ�kB��P�T=COZ*���cy�$��D*q6j�9=P9���W:6�I�Y���[S9�+��2�����w�_se�����) S���G���iq�-�e�?�I��/dNw�[V���̓���E�׺��ֽ�%��!	�'��"ݴ3,�~�K�^��P@���i� �r�M�Nr��(�5O z/���Ĩ�svW㰸�/�5jD������v������� gVÕ�Oo���'^ep�/��LV� ����$s;���3;Y֩Q��z��\�t>�>d�vC�J�͓i'�l��i?G|�ٯ]�K����唩Q�=�>s+L's�[U;L����\�m(q��|��/1�P\Ay4u��w�c�'ս���2^��c�d�(T����c���0ǽ}��~���	�/"��l��t}���)#�6�⟿�����6I�{�,tRz8���~�T]�|^��Gβ�fU�d���2���D�ܲ���* &<�� �E��D��v�\���ߘ�\���ʅ�� �Y�q��O��p>���L�L�~�h�����[�m��r�� H�-w-/�@-~�,��"hÃ��C�5�:��GҢ��¿�D�>��Td�A�ޥ�/�Y֎���/�[D������z5�1�6�;d�akҚ���_�h������e{��Y�_��RJ�Xd�B~CיÊT�Iy���4�1�? 
6�{����C_6ޛ	}���._�]B%����I����j�P@��D�Ko� q�o8[�hj;��8��_US�4Ek8o���S-�wݩ	g�����X��[�o-��jy��>:���u"mM �F^�gzbPJ_A�a�F%��j�{86g�͠H�?����  ��`�#�nf�$�q*u��#��2��H3�v�u:u��(#��خ�͑�p�����'�5y�n8sO�W��˝Cʉ,��%6\�W��,��o��ϱaW499�#+��k�o@���s{}H!��7�' dɇ����� !_k��F�K��g�=���U�O�ߍ��Q<���`���A����G���������������iZf�&h�.Q��0�Ô̘�>�h�p�y�c��ĸ��?����ddҝ۳�'k�}1�W����Lǁ�#Z�Ag�7ܤ��k��3oV&�ռ𫙉������&}[|)O��E���Ql���=�J`��[/]Xe���,�lK���5&�K�R�0���L�0S���y8��c%'��D9���N,���ޯ(���Z+C�bD����?,�H� P<w�eE5w��[F�ب�Ú�]�o��z�+�~�tr�T�ҭ?��I�̎u�ĥ9c`�]E�-k��� h���\�
�TGaYY�򗙺�_U�e��ޅ�,�@\_�.��գ�7�S�-Ee�(ߚT��R�b�i�K?"K��W�a}55dߐ�}�lv��+*�m��������������q��*�8�?:6�o�nWm�@sq�$-	��q((��Q2���p�%_�d��p��7��ѳ\�Cj��̆�
9�,���@nz]�+�BB�l'`AM�Ʌ�P�����?��h㍞��� Ӻ{��aDy�֍�h[�ڑ�FJ9{x��Ƥ��^3Ƶ-ٚ����g�=-��(�*�՗s����!�Y8J�u;0����;t�B�AD���z���\el4M�R���ws�T{_�B��S��,�����sm/&g_�l6�߿[���#�v�U+���������+�tnZ���g粄*u�0���ԑ@as��>*ʸ1�[��j�Z�u1y�W!��\u&iZ�z�ش_�]\Ɨ���M �Gsr��i�����(b�zt��6��W"��x[�yݺ�fی'��Y�2�'�ل}�At�_��y=�k��U��T+�/�޹��¹ȳ5*���@�B:e���f	�%��\9(��N���T���
�#�m���*�Kf�I;�;,.�����%�Ⱥrd)�C����ϛW	���L�h6vfU44��A>������������/��n7�$�4�8�#u��(P�םn��CۢA���H�Z���n�t.�
C~���<TC�G���b���ir+�x�
'̓\t3��"�����4	2��x��q���ك�I���+4�P�櫐��ݫ�T�b��I���^z�in���F��I���b��������	}%.�}��M��E['A�}�3���*��t�a�)-�#�x�gu�A�[�I�|�����yxr*�/i��{
y��d�`͓>��Y�cx��$�.��ع���l�n���<�3p8� {4�	)\�v[6A`,��M-�{<+���ͺx���᠈����״�P.?��!�RT��~"�L֥����4֫�76��� !��z�&�4�B��"��;�L�� ]J&v9dۢdy��S˱�B�	'�7���i�����*�.\�n �-�o-H�R�|�BQ\q(���k!\Z�ъ�S�/sQ��x��ְė�����$ܳ���"g(�\�QXi{���L?Q�{ԌBD��oD�@L�W�ќ�5g4��)xNU��f�83��&����Mن��.�n�H����$��:6�u0e������K��f��7�'�ǩ{U�B����]�1f��e��9h�LX�uV�~N���h|d��ӒfU�T0�g%}�3���:��뀻:Q����u�M���2oX�"wX���2Z���_��������P̛v�2�I �P�`�*[���%�Vi��T��f�P8�a���V8���jM!�;mȝ7=�����Q���)7�,��x�n1*6b *4�U/�\�P����l�U��s4�
�-�R���b�#ACWz;���r��}���6��Z�$�υ2�:3��nq�����X�t��+n2p��"�ʆ�AN}6��,B��;��uC� �ՇO��UK����,�ػ����ǐY�+?��k���JY��l �_�ؾ�X�9
��s�X��p�u6�K`�-hF+�̷c����#��1$�J<�/Z��u�6X$�����h|�ɼ'j>p∶���W�^�ךS���y_�������~E)�U�U
q���|~g6,��������ۺi쁼-S��V���O����~q�h��e����Τ�)b��6@�$[�����7�0���ȹ $�>����losѺ�G���dڗ��"5��[��Y(Ʀ\�	��*�g�>���@:s.�F�.YO�)��\B���l(��.���h>�]����k��I;࿧����yM�^9;�� I�~�}h�<ᦑ�II1{�JFO?7�|�m[:�
�F�K��o*�'�Yu���4_�N��2���V�b�6Bu�:5F�l��b��jU�m�5�S�58�,��JJa�Ķ�Mސ3���e}������}��:�/�59�O߫p�O���gSH��z�U1qk0$�	�9K7�ݞ��Hm��kt���r���߶8�b/����y9���?P>|)		���%d�(�Ju��ɵ{����� "�}ū��^k�y��k��N����]f
; Y�`݉�+�{w�7E$��t$i7֚n�Ul&��|��dK�f:]k^�fsq��9h��L����o�{4bB*b5'k%�����g�؜yG�r���"�a�+3����s)��C]���)m�q�:������]|M͚mk�HsH�o~�}'(��(�W���1�E��,*�	왹wwDJc��r��Ln�ua�#*�<cA�m��g�W�qF��/��r}&��p$��0���?��
���tc ݳ~N����,���z�DX�u��r��<��H�h��7����9��{��¹�Tj<S����[)?0��Z2s�J�F!2i��� BD��0?at�+�%z�Lc�{����0iF{�N�)��KM_�[��aj���7k��YV�� ���w�� Z"9��$���1{�.?� N�f�{|����U��?8����~�"��`::	���*L�<kŜ,����rC�)���K��F�������zؼU��'b����˚�W�$��A�y��k?�Q�pX�O�(0����r������!�l��K͹�&!UvT6�w4�M!߁�Έ�@LJZ���Y���G3�c����D�h;�秲��-�N�ݿ���>3�YA�4e!Ie�n��*��T��p����2,�B�yξZ���"��'\��Kz����m��'k��j��G �z[[C��Z5>U�D�-�&,e:�nk9��+	3IƵ0E��%��>L]��m��3Қ�3z���UXkUU�B�x�s, Z�B���%��F�j���)[z*h�'pd�)��5;;�|�����{���cI��cA~.?j�nAOU���i��퇛��6�k����&i�cfIJn�q�7�ڶ�r>����0�۔}��"�n���$�dD9�*Fl�>�1ׯ�i�F�a���zK������N��8Z���T������v㒖Rd��>/��9r�;���ТQ����$a|�<�-G�v�J؉EM�@�]���2Aa¥4��?A�k[.��R݅�_�	h�j`���ʳ��2��Xvd��+/�y��s;"%�ϣr���ɪ�vJ�u�WG�<��蝘����'{D/s��Ԙ���Q������0;{���+�!\T �R8���md|w�t��H��4^��h1_� �����]����L�k�6}:�S��yc��<�C%"-�'�xC�Q�-�D�w��>�2�ET>"ž��c�ڡI>�g��E01�Q_�/��Ը�+J�s�r�s#��v��������J�$�ҊB����=�ؒ�������4|�G������%�oh\c$+Ă�ā5�)����Ҵ�s�$]I�~�:��i��rqj���uu�}�w(�q̧T�T�E�.)iZM�O��L��/�k0�%���q�k~lg���=L�r��l/��	�2�9�5a�*>B����>n���ݙ!q=��
u�gG �:h���T�ٿI:�"^B�r[lZ��yY���A�Ni�!Iկ����.D�/����\�Zl�n��A6 ���C�F�ՠ�)6�V7�Q5;Rm�N?�*P�F���	ࡑ�$�B�ccK�ׇk�<o3�4zΆ��{7pks�0����<}��%�J]y�5L�H&����4��G�e�{n����x�O��S�8�A���|�fI��i��h�FB��y�l��"��2ĥ_��:�v�D�����ٺ�d�f*#7=��z�&�ϱ��&�pU���b'��P��+�$m�^J5LZ�U��g"b�e�_uq�U~�$�z��L��܉����efmU� ((��e^���3�d�������F���/L��y��M�0��XNM�JpH�m2��r_���� �l�@ .#�9>,��朋od��L`5^���<n&#�-�0f�?g�QD�W��'Uiq�]ng;>��3R���$�*���sRN�>~��Pb�~ �X�d�Ǘ�3� |��P6�;_w��
��gh�2{���ʱm;	�07���^�QT�}Կo5�J
K����d�+*b]��_6q;P8@��Ԋt�� XQ�C�s��-�^�y�������⠮��e�u��1s?�����=
�G;Q9T��_�8$3�g�&���S����H9�~��2��ȹ��:g�F�u��&xe����D�S�0s������yDݺ�_���DO�p�̺!� ���>��.�ƅ���?�8�Cj?p�	��l�x��#p��"�I�*��#{���㚶i�\OI�4���5��HtoQ�齧T܁��l���G�jh)�ض|}�.m(�DGhCSL�<H`�i~)il-x8�!}Ln��К�,����bDn���Ǎ$�����E�3Mv��k?WT���W]�ƛ����+����L.d���dL��2�*Xt  �1^����Uë2��%?�hi�O"�S>�IC������ُxk�A>��3��FC�
�?�LTh;���E�����8��zQHd�������>y
FVi� b�-�z�����u����u�ҙ���V3B�H�a$����>Qv��Z��K���k�=J׮��|NtV-�=���䚩�Y �%���О���-H�X��u%�|./``�"�t�k�,KU�6���j��k�c#$I��d� g�V����
Ǡ�a�\�TE�>���}Ʒ
�c�� �3�5洞.㻤g��Z|���ٱ6i"�-�1*�9�OBE��pv��]�}^zr��Ws�W k���j�q��T��3����k�9P�d��_[T�!:�DQ�Jt���Ⱦ��t͞w�>HJD�0�ѰN�V�y�)?Zw�$��v>��w�_��A�ɗ��|��CF�"ދ!Z� �XbW��A��T���
�מ�4�v#m�[�@/H��B��Q�X�W}���u;��_/��X�/���ק'��w��nT�!,C�	�����n[C@��)^
�@8�|�:">Z�hR~�����Cce�Wz&(7��տ�Y�! 
��A�y2I�oK#�jZ��D��B��Ŭ��+lT���e�;��c�u���Y�M��̨{k����N�o����\4�=FE��v�Jh+��dW�K!��7�� �6�p=(}2!}p-Uꌆ�)k-gW�k$
�.����ZȲg�{eA$�V�"�C����U���ŏ�&���n���>A�aNY��79�{���I������	�%6�V�"ei��&;��tR9�����`�$�T{:��M��{"��dT��܊����xC ����!�I%{2Ov�(�h<M��?��m��������8�|��?ݿ��b@������@tek:��H�"8�`��;����t*- � q�O��R�]��[wY˥.��r�F��aW	�ߞ��������y�G�븏��8Ϸ��lF�R��_��%e��m֞��n?R���	��ۤ�N�.Z���G{U������dGL��F��Z�˶bq^w����8��(�(?���"x�>m��<�m����^����2"H\>�� G�o�~_ҎD�l�cq��C���X�ǔ�&Wš�~�pںUbF�=�-~�����j
��@k%���B-��w��7��pVQc�%$x���>G�{�
{[eJh����3��tZ(E���-NT��"��B(�&�ȟp���|�:3��y�+���w��8Q��\h6s٬n��}���?�wׇc�E+�)�}��f�V2��&�v��'8�;��5���\���O���Oȣ�;,����,{Цa��T ��+�%���]g�W��tqPk~-h]�R}@?T8��s�q@�&�1;R�_i0�WE�+I�'4{f��`j����3I�M�|�A^�T�#1��0���x\�`jB��欶v)�ª݁��)��� �!�u�3���OЩ�??�C���'�B��Se���R��i��Q�J��'�Ouh�u߷':�Wl����|��t�a�Z�j���ڄ�#�2�|��Z��?*.9�����kN5�\��NyQsY�=��:�֦��)�d��=N�'n'�FW'ODp|����D���͈��B�'lR�x�rX�h��q�k68�*���b�"E��x���$Z�8iZ�.n=N���wY��"��Gz��p�Mr4&��֝(�wd���E�;j��>B�_P�/����_�=[��}��Q/$�����{$��y^v�u]�3ȳ��B:�Z`G�.|�̮~���xa��W||�ut�ڮ��
��m��@�736�\���߈��%J������%����ǳA;{+ղȈS��f�Pj���]
�Ӎ�T�110X&�f~�_��[AO�GḺ5�l8욋1����݃W'���s��^��d�����N(�,�:�=�E��Ξ��ZS���!' @��)��kVU��u���P�˲W�?�:�S�l<�����'SPS�H^��_L��GTG��14��7(p�	�a_@���x�/�,�8��#����E�l����u��ݥS�ޫǄ�B68��=H�茅�9;�M��s��l� �3�6�yw{p�����$�����-��(`�<��9�Ah3BT�͗8�]��(�;+:�6G�bc��5��uQ�bw�F�]����o�B1T48:�Mݯ�
GT-�{�����#?�̲�Gخ���Q��VK�a ����a��|M/E��dZt7����jZ�db/��xD�b�H��2�K�5����xFK��1���^��3����W�-������Y���?�LC_Ƃ�]鑸=rhR:��bl��3�I��ֲD���Je= �.]�� ����Ɋe�=�bc��K����8 �;�+`.��)�Ō+`���k��l��d�C�4�7!u�BٔB��،~M����c��{Q�q��ES(9�2�-���:gZ�א��6x7���M�����ޞ|>ї�e��ƴ�j� �������������I!ِ�Wl#7��-��]��
zRhK���8˔�}�Ƭ�!fBا���X<����YD�b[+���^z�����5�G}�'�L�"@y�t2���و��CO|�,ai$Ag �yR��r�����|��Y"�?�M�WlX�<�<�<es�ڛ׏ӟ�U��H��]�(;�yR��_�SL�oQ�������(A�tYQP�tH���d�82^�'_�4�i��]�=�sc�F���[�����(�
F��
eDMF�׉���L\do����k5�A�� ��s��Xz�_Y@��o^</�7w���E���՟�sހձ t=�r���՛^y�htܨ"Q�b^@�KDq�+�baO�����_��mLW�	!#K�c9�4��ZئK���P 9����G;�/�D0�+ŧj��yN�b�*�Y+��s Vf�1��_+Mk��lI�*�Cnʏu>�[�}�����i��;yҪ}��`���hM���E����s�]�9�q�d��x�5(���Pҷ�V��}�B���ܻ��?}ŜO͂`�R��?��v����R=U���cH'U_�g���l� \
���/98S�K���-�D:��{�]gI�7;�Ì��1��88�tN!0ߥx=��.�ZZ7��׾v¡w�SU8hn��[r���<�˺���z7gJ�E����s���~Z��#D<a��J�hS9��|"ZI�%D�)rq����jiu]&5��$OJ���p15�S�rg4��5�rMi��J�����S*��	�i
v�~1����n��凷���?K[T�zA�q�=��Qcm�%�
a?�ԫ�(�=��{�"�V$Ja��u��O�H�.�P3�R�$���%�3�K1N��
I���k_V$�8�N��qa�j��z�{n���Y�4������e�����؀�
jV���m��!˶$���B[X#%ډH?Th��Й�݄���еt���N���\t��r�_|(�M>�#����D�٢�����F���$_�ß>%��/�]��h�q_�5��`p��9��Ɛ/&�Z���q9 ��^��>�7�9�J��ҷ^e>.S���|�������~�~�J�z�4}t�%Ms����	T؟xYs�?~�w8��C�E&�Y�\�XlxVHYEB    ca58    2230��~������@E{�+��^w�<Y'�9;��[L�y}�U�����:�GP�<�C}Y �]��W�����\2��]��}�������h�@B�X���c���d�Q4����	�i��"������d�&���(X�~etcS0���%��F44�(?��Gtk�B�9��3�h�O��mx3_,߭�h����o�6W�#���l�)����'0�T_�Q�
�lT��C{��u�h"�U�@���<V
3�w���v��@DQ�g���U�+{��Ff"2ܪ�|�M��^e���6d�7�ޕ�C�OD̝�	��^��9�jv�0��''�4�CP�M��Pɸ�D�z ���ړ��/��N1Q��v\����s	���s��m��$f��oEn��-)���F7d�����cñbL���A��cB7�WVOV�I���6�k���Q�8���F j<�,�[��1�A1�~|���yu���u�����Q��L!P�DK���ve�X~�&.�Y��&
9�V�imm����F�umQp-�Gy�MM�;���#gO�B1m�²��ܟ,`�0[u����<��r���K��&s:�^w�b���*����!�x
�ɔ�i�
~b5��j�޳Q�Dk��BI�ڀ�Jp�߶~U�����.0�}�y���b���I`3UNv�}���?��l�3c�F��S\�RI�ko�v |L�!Y�k�t��rrJ�qg��Q�]�E�z��3Ct�".��Z�t�"�a��pp��M֜���&XYs�f6:��$~�%��tF�B��Φ����{���w��bb�G��1��{X��&��f�^Ĳl��A�a���Ϝ���l�$ha���F9��N�� N��/�z��8�,�:z�$��So����zW-uhtr�e�#<<�݃�U)"�V�:��4�?���C�M>ט���0@c�7���P��#���W�W�6��~�P
q��{���ð��p���u\-�y�����SF�'� ��"V����Yq#׆�	�؁Ψ�2�v���1�
bPm8DI��Ж���(�! �U.Ʊ3 �壹��!��Q>X�r�<]/?C�A�Nץl	a䴣��L,����ǝ�Ua�a��2���!P��
aЀ�p�W�6�E�e��瑳��#�|GqQ�ޅ4�[e�7���d��\���"t���H���,?/	���J�w���)x���@��"FR�!�����N��(���ٸk��|�ց��҂�-�iyL~u{��p�J��Y+[�o���g񞪉`��v����C�B�d#�T�C�����g�N:��������{�ａ�O|!=����}��2�8���, C;��[
��d
�j���Z�l砊v/� ��}�HwsǇ}�'����'B��UG�=q� 1%$��b�/�v&�����(ч�ǌ˧}��ku��U��g������=d�PC>��Ɵ�0ϥ�:���Q��ߛ�%��X4ǒ��%mZ��M� �S��-��<�S#vױ_��R4�{�<�c�Xmc��I��QT����!����\�P<�,�k�/H�ږ��,��I���S��S+�Q@�F�7����P�%0b�[zg
͐ث�;*��0�z]�ֺ�+�� _8�Ve?�.>9������D������I�6���M�g� ���~��0�j��7gP4�8}pT�G:�o�oX7��u�g &*,��Nq��~k���	�*} 0�8�&%����^p�\��s� ���BL��B?(;�e��`&V����qG#{x�A�/ً������71X�\k�CA[X���V��l�����l���J�����'�#�o,���>"�A'�+V#@��݅$�{��)>���Zc�huh"�5/� �5!�;����a�%2���9�t���G��Ʊ��B�Io�pgH5��4���fЬ�#Hv;�܌=���Åo��vs�il���wˡ>`N;��;뵦U�%l��XaE+�y�Մwѫ�1WGX`�	EA�-��X�
��"��� {ٜ�,�+��^/B��
!�'{�ZuA���*�܋6_k�K�cf��E=h�Ø��;�n�]N��Ju�~�y�!�	=(V��/ܣ!����*���b�w-黨���ٶE$P�T�W�0Rv;x�֜���\��b�R�V���V�#��Z �y"���h�XzԵ�-U
Qm-�L'�CO��
62������D������iֶX�]� T%��qW~P�]� ڭcu��,��<�w���Q�їc@�C��W;g7�E7XA�+�Ө\�uw����g��<?:�����㴪;��������~J@�K<v�)�`�k�?�M�FGw���F��ʙ���q�5K���g���$�C������Pg6��˟깁f��۽�1`u�����r ��������j' ��q`�����cZR�\���pcؔ�@�Bĺ��W9�ZW�[���gSf3I�>>���	��&���8sܤW��լ'�^�s���}��S��,��iv�7�p�j]���c����s���pN��k,l�wwU��; ���<5� d�-��R1�3�$��%������#�Aͻ�t@}۸���Ԉ�ʄ[��g��+nf7/���D������LӬ%5��a�adk������WG�E��k!]��ڨ�
��&^�j�ߝ&x���#�
��p�u�>i�<M����;��><�ӕx�.B�U�P��#�r@�{����4S=�`9w��0:�#VD��,n��a ]̋�DeK"U���V��9:����兒WգR}{
c�hǾM��QWB͒�����X�6ͤ���c�v�@j����(1^���W��G�� Qmu��hfZ9�T�Yh�����6h*�w�Ƶ�K[��;�`ڜ��h}������1�M(��Y�:��[�����֒���pU�{�",���-6�=�?nx���0xb�հ�Kd��$d��%�n��n[t�j�8lE����!B&��(n�g�?���
���F����-T�=c���J����פo�0A?t�	_�Q>�!^L��������~��e|s���#���h+]��G��(RE�v7!��h��Ar&�^"r��1�b�e��d�y"��5�l�����PW�^��t�v[�,:98ON��W�Z&��F�͊�S���D�:�w�1$�+pg2F�������&,�}�Q��a��iBsb�!*�aO�?��q��▪y-��!�������Z�|&{��h;8��I	j&��ɴ����T!*׹H�.�6/h�[��t-�1$tLO(��iR�g�'��@k�� @��`�D����eǽ0@�a�&�-�5�r���}l�ܻ�:ZC;�"[��ab���t���U=.�m\_R������:.�p :����S#I�1>�[ǫ]}�`E��_K�B"^�/uy>b���$��*.��g-��N\�Z �WjkO�c���Q�� �� "�FK����,>��_��U��>�2NQ�c׬<�<sLN�\�"!��:s���� g츛פ���v���On����}�'#��
z�����sEL0���+���RQ�C�aq�FFc�T�1X�9�V�gO��.�y@-u����FI>�	W�c�F��bͥ���j�A#%���Wj�O"����t���j�š��"�C�DDg/�[\�*M8V����:�8I؛�ʇ_J��?x�9C"���r��JN
��5~8id5�T�r7 ���o���;r;T��GO�OIW��IU��/����Ϥ&��qU҇6��84ƹ�ph�fCޥ�m�f���Te�LX&"�mx�Z��G�P`:�	vZ����Ϊ�%�"�uCWƻu���
~6�jg�&Ð����о��%L����GQ��%JV�M�[�;�kѽ��� �y�aoZ��є��G�5ۉ���"�������8�z�����\q8���˓*��l��| c��<Ϩ�u3*G�Y�ۂ���A���
KC�V�7�a�RqG,M�ߴ�P��}�+����c�/�~�!u&ĬZ�]�C��<K����4(�����Q����J�J{LPpcr5��c�{d��ñ0��^��aN��+
j.�U�d����y��d6i���zI�6�@'pOc��x����V�3��E)t�����9�N$1?��A�<��H���MO�=ϋ��s��Nd���Mm`���
�q�\8��t�/L(����֍�`�z��H�r�I,7(e�<�7��toa�]k�@���{�,��(��������$ҿF�I�F��\�t��-�)=,��8�����oF����l6N� ��	���]PA��o��B;�.,P��jx�z_�r��k�����eH�8�ϲ�Q�>HB�7���"�GF1��"�U�V�FTT�H˗4gt���}orb��������35�*դ�NO���PӞ(�)�pЦJt� JS���s��c�ԡhW��d�1s;�1A9�D��2V|J�Мh�un�[��֧�6��I6�8�"��z�G5�lt�{�Jw��h�ٮ��8���DЁ~<����Vzś*p���Ɋ8��!��J���� ���ajքD-����WVd3;�� T�$��� K*��b��!vW��b�H�_"��^�gr���T<!<�+X�G-އ����Lق�MC�0[w<dUj����c��E���Y����4�-{��R���Sg?���|�I�ֺ��V⭙:1���?We�"}^�~��E����2{�6����C��$�Y�bV��S�R��!'i`)B�9�����8��S4�/�
�Z0��_�6�5u��S�)*к7Ĝ�M��%'c��S)�2�>�;҉ڐ�<Ӕ)�S�#H}p�Q^���<���Y -/��M��ܢL8>�%�*?�߶�_���`v��K#���+��@o(!�]xP����R�?���C��������z�����s{�<W�	�'�3i��f]�f������xpнF!)?����� K�2��5X��s��
K�x��A�mm������T�v��_��.�c�z��"�m��в�r�Z0O�%ߠeRqgc�`[<%��o�'��!�;�'�����3�.��:�D�LV��c%ۉ��i#&rp�7sU�j�G'`@l��|o��z򰐁дFce*rv�D}}M�N0���l9>�U"i��"�MB+���=w���^�*�7EK�����9��OJ%J�B$W��
��-�������~n��.b9��m��@�p��u�nq̺��f,R�ϏT.�b8�C�9�i�!
�(ݟj�]�~�\w��Bp]���nY蝍����.��d�Cp�͌Yd(�:=yo���Nש�pa$�3t}���#>�Q�2)Tio,�'+@긁F�f�{�G3��P��\u�)�=1��dm���aH����V��(���z�	a��b���g�`'�Ø�/��:��:d����Y��0��p���'�+G�y��4����30wp���1��<�W�����#ҋ[��?�'f�,�jp%�,���V場 �N�ř0�+7N&��Mέ}��o���ω3�r޼�WI��w���*�!%\��U�&����1��	�o
λ�/�*�,'��r+����x�*���T���)��,m2z��~��_�ھ�4~�| �:2����v�*}��WX�0  �	��I��4�pE42��oyA��~�hmByBV5��͍>̛s�����J�ۊ� hL R�����ڲ"1h��5	^��f�f�)�{w�`^@������}\���0WEs6R��� �
���V�
��%;�qqvp{�ZVP��3�)N�Bt�h�ad��s���/�;�eL�(��PJw}xUE�iֽ�p���n52o^�����ǨM{��`�z�Upr��J�lNQU��-�%��6���c%,2"H�����s�l�mf�Z����D#�AiH�@	��6���tu�<�5�3��.�j�](#s����^2�Z���<�ނ�&21��>=x��w�0���\�[�h�4%�/��F$�r�pS�s�7o���KILBVn�m�F�Ṻ�i��)H�,/1��������="�w�λP,��{���`��rţQ�����K��[�3�?�1��ޛ���"�� ����Z��`\�r^ �ڧ�ivi���5���Y����� �cY֛%ee�����~�J���@���A���.j�j!�����D����,�&��L�-�@�B�U⿞j ��=*
#������"�(]���O8��:X��l�Q"�<^��r[�	#?bN��:6Y����U������VY��rٿ�mN��N��e��ql��cIz5���k�����6�A�z�=�
�����r.��`(A�����Ey��"���8�K�p�:�-͘���wY1�|�ޗ��#�%ly�'�+����>�2����]��A�Q9������ZN6�Xq]�����Ǧ�fRZ2=!X��
��e���ԙx�����BE5�lS���j6q�x��!`��̎���~�&�6Bm��*�6P����f?�J��It��,~?.�0t�?+Km�!�E���o8Z&��)(�S����T�U�M߻Y�,�ᠭ����y������P��h����K{���p&�;���?�[�Wl	ςO�RlhO��F�=��݋W/pC��K�5ܤ`�v�T�3Mp7Pg��+�o|Y����Yڃn��u��� Б[�#�����ȹ��g�N=��޸1���9gf����f�䏒\�P�Zr��g�}���ѳ(�+�@ �Ǉ-Cp]�%��$����|��SX����/�i�������= &ڤ��E"��?�~`��MJ(�� �0���O0������]_0�{��D����YN���N�DMu�Ͽ�I�RB2i���j�,e�+4�.����bO]sGuh��
��E�cA���?@����O��?�N����&�>ٌ�1�&S
�QGr
MF�Mi��\�,�3����@%�À���vHLuɞ�P10uO�^gg��N�G]�ҹF5	����=O�2*��T�
"��GK�*I�_!�λ96X�CPs��e�ҰL���u�o�:���J�n�������1���{,ݣ��-�MŵZv.��R���
�)k �����w�K��)�N��k�[x�`�tG��qP�>�n��D�Z-�M�rod�4�F��m�� z;������s7��nlh5+�4��f��L�֭��1Ά���)� <&�.OĨ�w��u�2�X@�a'3xp����N�2O�I��wV�2���sö�
��D �#�< �
�[�$��:��M{�놌mu�-�bdSy4�<�$�K����Z'����fpiI���~�Hk�WU)=���+��k���Y0:c�ߝ��
����i�
�=A��k'���*��Ǧ���c�n�_C�����:�X �
��!\�^_�L^'���T�"`6;4�YK�j䗾E+�S)�d���Lc��Pl����1��%�4C<�!ٻv�r"��ÿ3b��}�X��;��;�������<�md�>c�Sz[�U �p�aƝ3���#����hpq��:-���5��s�;�efì�[��,��I�V�@ir��!a��laN+,i	Q06�Y�q�PM�`4���z?w\�7�~U��M�w�<���4To�0`�W&n�d�p
�O�F�ch'���w�Z���Ⱥ��\O|�T{�/]n��cx��wZ�Q�%2�x�b\��d%��AeHM��cm�Y"���E�e���P B�g1[�+N��(�������4t]=�k��������n���D���t��+���*P����R��"�	��Y�D�=�rHƭ�ر�sO�]��%���b'8h�"���k�D���;�d�5��2���gK��9$��)�� �rX�&�.�ڛ3��y5�"�Ѫ�`�Y�Z6_��(�հbnR$&�6T��J��� Ň��킸� ~(]7p=%�� �ݚ��#�Is�c���1�6�!�b��8��
ټ/H|�aȵO|�wRV�T����������IΔ+��-8W��V�-;����4GB�By^��]d�U|P�Sʭ7�!�@n�b�J��Iν:��j�֭	m��A8�yz��<6���u�~"Ac]D�^*T�j4o,!X�E~>�V�Y��L��P��r{8�f��Vm1�X_�a�d���)T����w�����d>;��\��Z$��l}� ��0lND�RI��bh�	�:6UT��?���1b��������>��������lq�F���~�l�*���f+�@��(�U"0�c	�Nl5�S���q����������f��m���t/�������1G��Z�Z���������(���D e��=�7�V�yZ}����r�������P�\�m"Ӳ<�b���I.�>�&��%^[�-V$3sҡ2�6r��N���2�c�4@