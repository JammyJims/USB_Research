XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&��{N}�������+<\�Ȅ��(`}���o-��]1� fL4pM�R"���t�Q
�aM,0��e۔T����P��u�QoM4��Y�I����v�U���F2XI�/����Ct�,V�,�@��X�д��K��[
�>X)l��!�W�D�n�By~�A�7��_Z�u�^�2o�/�A���T�����v*��L;�p!��!g4���hM�~��t��M+t� �D]]&gQ�i�����e��ϓ�?y�?����
�v|�iȢ�?�?���-�>Sj�p��C>�U��Ux<;��T� z9�Ծ������I]W����l��_�>�Lǃ2aa(��1�U�!doFm�&/<|4���9��!�;���9qS����	�)lZ�6/S�X��O�I�)r���G���B
bj���S�Q���f�kF��㳴ϥ�1���,���K�ÖD�=>B���&��2h���*��z\m��S��ICy�1����L�X[��݂����#���� �O�r�uj"㭕�2�Dά-�is�bs���֨�w���b]��P�g�����K����s�����E���C�K�o��ް*�� NU3���
�UwTz��Ē�>��^�msTd�m,^�}
}�U�r��<��5��X.�tT3�2M��-8���H��TO���smh2s�x�p�KÉ"]��̶����3#��Akֻ>[[�vj�+�C�߰Ӊ,��iXlxVHYEB    2580     bd0]e�so��߶���~h��� �]�g�!Αʸ4E���;��v���߂�� +�n�T:��g�2ص%2���ms���,~H��э�A�v|�Him�\m�=�����C�2c���aP` $sLtL3�6agL��.�c6<rI	��}�힭�~����%8��ߕ��&��f���2U"݆����?MT�s8c��V�e���.�|�{�0�SE6ƕ���ޤB-�D��2Y���0q�O)����)�ԥ��?= `*�چQ`��.��y���9�p��o Nd�"֢q`�ꉵ�p/6\��� �4\���@Y�z�>@��mb5���it`���*�-�<=N\ 驵��;��Z�]��p0�]�om�Tm��9�S���w�K�BHwnZ��+�������u"X�zO�椡"Q�Ό�uw�6*si�:'�I�W���[��_`��"Pb�p<j�>xz	��Գ*i�����ؠ��Xl��mh�$M����z\�q���f݆�6�����ٽ�T$�R����1�%�+$�{9��vo��Y^qy�C �rV4��G�5�n�:s�j"\�-�
S/sIQ��N�T��o�H=��nZ+�AM�R��zgH���<�֎����-���k4	�f.">�I�t����Z}�g����t źc��
���<�53rt
��x�9+�|2��2�l��)��Jf���x����ޥ�I?��w�X�T®�Y���â�zNO(9��j%Y��}�٢���� �'�F�9R��0���Q(;y�
5|�Y�Mj���Gk@��B)P��y'��R�椓Bh�q��FYRgB$uN�}�Q�א�SqN���W$�1��H��RU��Q:��X]��q�b��f���ˢ}Ѳ��~�~�V�|a�3���b�aǡ����aC�UD��A8j{�����q�A���{�R���8�
h�t�8\T�ILPjʝs��tTB�	����dc1���@�J�9@�(>�8�[��f�>�Ѫ6���8����A��:���ތ���7`^:Ք�`�}*Q*T���G��7<�:o��S��
�lb�����T�I�O��d��k:��H�Қ^�(ㄣ��vb5˘y�t���$�=LW�dM�_���'��1�d����p��� _�h�x�����SN v�"��c��	$D�&�	��-'���4�$ώ3��U���O����%^����Ĕ�]��
j�`]�J#k���
��OC�95 �W?�I.�.@���ä������#u���Ic��h���,t)���^�Ok��
�1�>fѫ��e+"?��a�6M�J\P��.�\f#��]@Ŗ�A�:�$) ��l���-X4�=$���3��"݆%n~�d{�o#Z�q�$H̛W�}�4A_�(��o؀'���T�D��ⅇ�'?�6 �u��������}�Pn���od@(4�#
S+"
Q?�+W�4<��WZB�0�x��N+4�ngf�w(��o�"M5�7�$-dѥ�cb8Q�^ �q�+����|�
��f��L�{s�G�a�m�+�A�ț�h~�H���WZ�i���A{��lS�!W��Z�B���,���� $΂�O�=����� �<���D����u��,f�[k����1#������C���CM����B��p�9в����*����"��F1��
u:�������'���`/��0.�%D2��܅�4nzW���V� ㏫Z�VZ�LV����h�2&R�Kd�ۉ�_��������m]H�oz8�=@j�N��-S���]N�@��4
�<��z}�Ee�i5�jl�$.:��8�v�s��1ȃ�S ��7B��Z��v��^��7��.�z��W�7��1)mK4�����̸QJ2��"&*�$eAYWI���8��ޠ� ����:�s�����������,���%!�ܫ�*�#�<_�Me�C���!`�Y��OeZ��;��n��:ui.AA%����~@oҁ��1	fm��JN�>��;���5�[�����?�|���3����݂B�ӡ��c��[�¾/&v�nژa�f�x�A���M!=K�Ʈ�_���:�=\2�����X׼�!C���0��u�� ��"�L���1���t�x�5������\��`���$;��>���	/��t,E������uv;8L�qAi�>�BXl)�w�b#ˋ�Tn �XYa��Z�u��>@�y��ZbՎӯ|q�6�O���4l�8Xڸ�Q�"g�NߒϐSb��'su��]�jX����Q|�03L��"��<�#����S<�*��� h�
o�@�",����<Q"����"ާ4靖?Cq��AOS������A5z�J�8�������Zz(�<�@�N�b�1���Y]�
|�¸$o^�_��l�F��~�iE��]���4�$����uh���k�d!by�+������Vy�;�y��6T��F�|�z��4�4x�� 2b1�~�B܎4�\�Tk��΢P�BR\P:2�VX�ua�����2\�5Nz�G�ʓ����T1��¹������Ǿ�S9)&]�:r6�e�P�hU�����T���{;����*���� e�������`ȝ!��+Zr�R� �Wl[�X�v� S�"���I�t��`�
��G��" f� #���J3�,i�z�ֵ:��DC��@�^wUB�;�۠�Y�!Ps|UfY��J�����>�@;Cђ$�cQ�Ћ/����ԑĕ����]Y����1�"WNx�}�A�������3xw��;��B��n�M��9_���u8�U)(1���.�׼Y-��#�iz&�+��)h�jtv��u�@��C ���=\�����1��UUu
�E��Ų����5�Ft-�Wm����VqV;8U�@��dl࣍S��4��������~_'z�Ә�a2��S˼#��0���q!���f�r/ܜ�x����=�2W��{l��P