XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����C�K���� /p��8���Q���#�.��zݑ:q�oc�@�x����P�O&��`4n{V���!e��ֳ��.'{4;.}RtqD^��1R�fͅ�+P��ԍ�|�u��>�k%��,���@���3wF�\��A��wj	��#x��`1�L��O*��s{6!���c��a�G�䦌`���\Q��A��Q�w��a�B��F�,<�DK諀phs��p�+ǲ���d��B��Viz������RB��&e2k�foQ��#q�m���u<��!���tw�/BB�����7ms3%M��a1@.ۚ��}>��� �j�_nq[����G��G]�̳�z�]�=���nHa�*�x������
1��πG/��	�T���ШsYC;���?hkAsu�;����/�o�,�RD�&,���#U�G�]�w��on4�`P��T.����X`S2,�#Z��s7�zJ'>���0c������*����J;��3Ց	X_��N�h��_�����G���I4�c�ve(����	+��2G��9{;T��������*י�����%�_C��:6d ,"�m �FvĒ��p�,����;�..6:&�Q��=���B��"S.��؏�Q���mB!#E�c��e<�/��~�nʒ["�����p�R��=��0nX�1c�ɘ]�[��\�`���0���S��!.*���=f�����M$R]\ؐE�-��]��cs�XlxVHYEB    641e    13c0�s2;����ֺ�ǡOi�?��<*���i�*��]p>�+������ӽ���X�y1���=Vn��I�5�-��X4� �^-a��i��]I>W0b0]�e�iL~o�O��xp(�Vm�O�����XH`Ze��V>��t=J��`r3Fm�/ä��'V��f���?`���D�����<#+�� �XYƈ_Q[�*�Ӡ�dDK�(M1�jS&���m�>��|��a]!�h)~Yyu�mm�Y凝�>� �ZC�p}�iNۡ;$y��-G�:��K���[����� (%Dc�`ՠnk��� |�����ۣ���!��Z�Ȕ���АG�/)0v�-R��(C�ٶ�&�P'�Nm>��V�Ŗ��_��hKyE��k���i�S��Pћ,��ɱcc�cL��N`����F!���`�1dƋa�:赲��FrH��Pr�ݏ��*��
�C��~�޳���\,�G��i���]_~�}��t"g�C�U�m���K�"R$οO�i>Mg��H�n��K�&���$O��a�j_�(�Ո	����6`ŹLm{�є���ޑ��Lh����?M���+�n'���ک��F(bF�N�-�+g%Nc�"�< ^#����9(�� �����̱�(���(K	��H��`�b��K�%1��Z��5�7F���O������j�Xh��zz �LױqZW���X��~�����D��S�R�r��4������OYb`#hLn��݉�ˍ��Þ��t;S�c:b���k���'��It�����ɏ���P��j1���Z���#��
I���-�c�[!�o�{N)�O�fƸ��@�g�]�ih�/Ț�/_C�4�@��t�t6n���,7��E���j2}'�o�[����:�1��^�:����\�{R��5m,�:J����b�	��wZ�S����;�E	t��f^�j� ��3'����f��b�6뉛��.?G�\��j�Uj�Ѹ՚'�&2�i^N޸���Q��b>�����x��RLiJK�m�.�y�qo#3���t(#��޵����̚na%��U�B}���8�|%�ߺW��Sq� ֨I��ݒ���N���W���m�]��PE��q^�#
��L��#_)��Ι5B'�Q�U[�%P�� �2�:��NC��k;�j�&:�_�����a�ց��5�)�x(�)|�/z�U���55T��<Ɗ��֋�_�b���0�M�O3�5�X����y�rg�ۓ���	��RI9���A�kM�m��i;/�9PH"Q�����>�DH/#����8�p�@;�Nx%���N���)�l�ٽ���;���^�o�86�_��ۣ�j�׵+R�:ĺ#����j D؂M����WY��8am.�z��v?��e_����>M' �SlHm�+$T=��㐼Z묳8vh}搒�
 64��.����R/�W��/ο�=�5m�l(#[�ҩ�� f����HG���wPanún�L�}�+R���utV��J
�v�y�2?y��$O��t@��Ǵ��,৵���˛,g!K`�_]l&,ն���ݣ�v�����r���*���L��Iެ��V��kR�T*��ِ;����]|��N��>���f�e2VV{V��.mnχ�2?��u�g#_ ���IvOy��8F�|��N�i����OQ9�e��ت7)�W��Cۂ�)�%�ʾ]p��r����uM�o�R.O��>����QX|��*�b<v{��y��p�2�ݵ�6�4��*�Z� D���Np���<��`��mO5�W�J�>�ps��
�1�TY�	+C?�#2��,Wj��#z��Q>�����~"]a�{�7����Mm�o^�Wo?��j&����H�]^p����)��@�j�MƬ�Q50Y+��
!�z[$�lHЩ.y&�Q��)I+��Rį��f��Gb������)��d[%�^� Љksr,����5o�ׁ�Tm����m�Avf��4Bk�N�\
����V�掋?[�a�>d3��w��Jg	��!|��K����p.�2��ag���^��2���d!L:T�Įv��*"	�Ӧ�]5T�e	,�?�R���uI���pW�k��\�����w��jg�ai��J�g��Ci@�p���	�n�d���T�|��}M�K	XIB��3IHk����V�'h��P���DQ1���qe.2�y>xRɐ��6�rr�=�$�ɈB��Ia��d�Eb�Hג5�<�Oj��C�.	�Ĺ����yr���a�pjVos���/�����I~�\�㷿�͍6�fgF-����٤M8�+ĈAj���4���o�ħ��C/1YN��o0��Ŋ��jV �(���
��|
q�#�Y���ߣf'��eX�O������� �X\�ln
U�n/������m�!Equ�KŻ&�{"��%���i�9��SJ�m��( "��$�A��g|�M�����IS'���-��W�1����D�Z�\�u
���Ǥ�%�tw�?N ���@{�����(�i�?��ֳ+-��ҧݱ�p�c[�i(�Ԝs��n����*G�gx���͆�L	�S9j���SŪ��Y�1)̀A�#�2�(��� �@H&�}1��K��m\Cx�(P>(����nح8�E:;�O���o�>�r�<S�qQN���`�C!�ٙm�;y�����@������!i
��";͡p��������,�5�����Շ�/�1�l�m
x�B�˕�r
�����$�����=ڒ�)�ǎf��%<�3�c�p������6��zȪb\@�
�O� ̆���v�	X��]n� i�9B���y�ŅM(�!�?Zm�������:�-&����n�l,m�5!�8:C3�=��������7����{zX�x��9�7u��'5�\^�[=�/S���U�K�{�ʯj�rFOc�e/*0"&�'�#���BFu�M��\�	���{�[���"��8����W��Z���G0N,�Gףw���sn2�!U*�R�V�QU�������;��C��"�ɜ��0�'��|�������͎��GA{ 
��N@�rT=q�?E�"�m��t����q��O�*ފ�_�R�/pA��N>WQצ��M9X�g9��6r��� ��O+�fXO�=���6o1���9��m�:e[W$�H(�g�&O����M�r�ǳ�?F=�Y�$*ed0OL�M3_]��5�����/ꌖ���H�Ė_!��(Rي���3Y���o�լ4��"�Kբ%�Hq�>�ɬNJ�G[�$��H�7�R�L%{�d_���KԷ�jTa7�P���QR<��ܐne`X�/��wݼ�t��K�5>�����Zzq�����'i~�]��%#����Jy����[��r�kdO�U��ILf!A;�>A����x�u�)�n�|������B\_����7�aɟ�� щW�d���D��^�
�٨*���M���As������5f*��+���}=�@�V�dV�ӳ��@ǫx�ll����F ي����[@9�q~�:�ʌ����i_�g�<P�����u�8�PH�Ư���˱��fq����ߜ,�y몧�����Ԍ��\��r#H?s�ם��
��~���g<�@����dm�o�x��u�l�J��k�X��' v؋�7�F<�'�p�]vr�}yAU�'%���٧=�/C��]:���O,�'�l1ʒ-)���֩e����c����ˑ>��Q��Zt�CU�w8({K�;b8���"%�j�������^۞�u��K��4�����<N�◚`c�|�h���x�q0�����C�;C����y�m�m�O�S�&lx%���H�0��4���Z�]�O�fĥ6���)!���G�l�����h1��~��"�4��*=%��4�2oNX��28�K�J�2���\����Av2�<��g�͜�K��?"-S&"��x�1��`� W���.~{�1��0���5N��z(�~R���T>��~_l���Z7U�`��7P�6�3�m1�vsl~�&��۪4�{whgҩA��9�V8g�f�������Pv��=�{���2[$.���-�Y��࡛
!cn(;���tK
%�A=�����>h�]�?]����j�]m��⛝i*[�������RY7V��"[r:�[;��%wd�7�%H���"0�sv��%X7�0�r����Kpww�x$��[G��/�!csGfwK�X�Y<0Hx�7��c��<�u��[�ђ�{�>�Ӭ�j��'��)�s�:^��lq��{�������S2Y<\�zNZ,��Ŋ*�2Pr�a�;�*$=/��揫�!�1|�	� f�/
�pf�喿�3,�A�?$�n/*ؐ�mk��S*�ﯠبd��;�����o�gڏ�a�S�zF���'Xi.�׵_N�X�fC��,Z$R�1�3��+A�	�� �]3�����o���[��(�xz��gw�Tq�!7^:��w8<S�9�1������U>~(�����xE%A�	�]�,2lJǚnN3�Ǣ���hG爮���ur�Q�h&K���:����������I��bkO��6��~��o,-L�4��z�{�"��J'eT
{�h�_mfx8�� �
c�Y1�b���&��SD.>7����&�V�� ٤�D���v��e��|��9�����?�GN����Y`��k+jTt~��l�'���t�
�M���'1N_�U��X�#�s��;�T/]���b������"Tz���6� �Q0U��H�HK>Ֆ��7�	{�>:�����=����>�K9V*�q2-M�ȷei����T��!� -t,ޕ9���^Z�`5�O[G�e�q����'�
auK4��{����aN!H����n^|