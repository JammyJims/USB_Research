XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�R�u�ު�7���C5y݂g�O��4���]-�ˆ� �.��6�[G2RQ��g!B��=\�p!����6+���|,H}��Jl���r��;p=�;*؍�]�e������犾_)����Y���Q-��#z��D<wM�|r im�	ᩤ$�H{7���D�F��BވL���e��ipIÇ:�X�~3H��ׇZ�ڭ�ai��Ŏ%�����	tD�_3�����2�����LN�`��ȣ�H>�{/{�Ko���4ݯ-�����J��2�P�E�|��e �L5�贬IyR�Ԕ��O)@Ԧy�W)�-	�@;;�#Qzu6r���p���tpr7K�>��Œ�}X�f�w����v%�,J^��ʞ(�h�e^h[�n��F9,�|q�J=�����em6��`��(Z�N��ؐ�ΘO߁"��(�3�_�F�G�j(��3o�Κ���qUu ���5@���ua����p���.��l�Q��1��`��y5�k�O�c�90��i��ґ��a�@���vN��+�Y0�X4
v�a�]Q:@,�vw��;���˔���{r�#M�6��~R�&~��"E�b)���r(Gۭφ�⢫w�]�}]��$�k����<��-z^]�3������*��|t =������Ǜ�rr�rj�U�����n$�0#�|\����[�'�#�L=������J8�k>���+V��9���o*/�y�9��+ʨ�DW1ZB_��y2�;�>�?iXlxVHYEB    fa00    1a90�VF?[Փ���2�N ,��^�����"�e�.��P.�F�֣�±dv��y���&ac�IVJ�2ܵ�7RMcu>N�9�����z�@4���)�,��GN`���L��@1�pڍ�G)�"�~�3R����c��˃^s�$$��ݘ�>b��;��?d%���5��Y�F����	*���Ǯg�e�V_��h� ���G��!��8��c�{7��P��M�?ջah�5�z�Խڍ�Ȫ�}]�^g�mğ�,��o�[�ʸ�eEI��I�Ǉ�2��BB(P�9�d!��6�)�(c� ��&��>"�0�0�o��e�s.]7����?S=��T��mOBݮ5	V�;]���W������ڗo�����*��Y����D��B�ޑ)dg����Q����5����ٖ�����B��B���	&+���y>K̳鐑lyW�9�ί@��w�9p��KX�dN�U��DX�ql��7��D��"jD�U��{�����|��A��z���ِ��2�0ԛ)x>��\��W��K��#��Fxe-t  ?"0�:�Wư�̏o0F3�L����eO~z�׋��v���B���p��Z@*�j�����q����;Q���_bgm�v��˯�'>��5<� �<���y*f���C��^�R��H>"z@�;�n���r��9��P&�B�~���gdb4Ps����8��f���D�x�ٱ����������A��a5�w��`t{67�,	I:�7�Pn*��F�(�/���nPȚ�L r�d��HD's�D�[P�&ߢg�X>0�L�?]�b�CijW�m#~k�L��B�ʝ��+ b�SL�0��K/���Z�0�6
;Q�ď��[�`�X��`�����ϾЀɰ�N��:4jMP�? �6,�fm#A��xfneX���Q�КI(A�y�w�!��\T0MA��ْh4xj>���A��ף��;h�>�	~���RV�A~�f9duo�zC�Q��5����{��[�XE�T��B�$���]�>`A �-���,�a�Xn�		�C��o��TG<^o��,>zh��P��'�xX�G��E��$R�\)ao�����R�?웂�T����ù� �Y���p`3=���2N�d���6:��'�8)���`�i��]���p��R�W4�f�!//�xF�� OKyr�d�U�NLJH���|���l�J$&�0�uBup\��Z)t��P�dɸ�__�C �vGҺ��h���Y)�i��X�t%{�ӯ�r��<�zbr�u��>�;nJE��$�������t!����Db�B��|&/>M��M�p�8P��ǵ�XbaX���.���Q6?D^l��d�<�ka����Y�J,�4��]��@�O�{�I��Wl9�+%h�ly�����'�=����R�� �&�J�LAnB�ă}��	�ٸ�¸h�eC� �y���� t�4dY�����R&��� ����[����,����lN^��xs����=b���Ie\�n�1[���*�$�jqs$��8��#�RsK�G�y��C��������k܈��4S=~��[	��n�SϺL�����k{˰掬� ��t��m���|`�k�>�~��F-������ /�e�̀Wi!T�l1�\�E��⺇�h�#l��C���W��;�:�)c��)t����!r��|QnQ���+��]b�{:��`��΃ǻ��Hd6����o�C5���m��ڦ |nԁzk��?L~@]س�
[�ϕ�dQ�i.�e��oS1mMzMf+���8�468�d�����w�&s�M���y��+�[��{i����0OT[��H\��S��U�r���~�u��C�^�U�򡬎��
��:�K�t _��A��ya��:\���q��Ϻ(�?F��F'\�!�Jc���K�;�3U��2vy��n�>P�<n)�����-���.�y���\|�W�v;�aӀ ICB(=I(8;#hF���� Fr��4M$�NȄ��fnk�����P��$�D�u�$*yK�_�@���ȏ�%C�>�P�m9R�F��8�yT��,G�w���V�rUv� e$��cF��_v������	M�a�Ld��:Ōd�
V�>��t�P���d�a-V���o�����=�i��u�ӳg�Y���_���W�G�V
|�ı��3���ʸ��Vi�����P��襚�׫��"���汏g]G�~�M&�_4n�Ů�m��Bk��s]Th?�z�ކ{e�'P���kl�3K1+T \͍zh�a��J��.��!9�෧�0da��B:ƅ?�ؙ�{�&�f��>��|�q;����[JA�T�Q�<���<ɛ�g���_����е�%C�Q�u��}v\{�.�*NC>��+5#�~V���\��H)J���>�� n��%�v�Ј�Hȶ�c$�|��H��� ���w����V�bD�R4���}��q��򁽇@*`73F�?]�΍��Ll6u�K�\�����1�m O7��	4a�u�uo��%��j�*ԏMک�1$�M[�\�ދl�r�G�~0�Ś�i���?ϊ%�Y޵�ĳ�	�ጎ��&{��R��X.F\�.
6��:ㄵ��UI��<�^+�a�gY�mRU��:�U�\r�'i�i+F�ܔ[X�^b��b�a�~;Q���Q闘�;G�Z(��zГ5�A�1�r'��7Vh��Gz=�>��#��D�;r�N��xD�����%��֔m|	n��J:���V�%Gw�&dfZ������}I_m�s�ڛ��CIjP>YU}m)�����(�fv7,8	��b�P%���iT���1P��L�/C��A�_���[�e�$
��A���hrsDv̄8|9�t��:��Mʍ��������RzFQ!���B=�u��:YP�u^$#9��<*~G�UE��Yc�i�t�J9#�8����w���W`"��V)��=�sτ�
@����Vf�9D���D+���>X�;�A"gJY7&~����O5S��? =���=��5ި����s�e��������gbM2݋�@�:/^�_!UH��b�n<�St_w��U�v�y�h�CA�O��d�J������O�q�J��M��a�C�ѽ�$z|�4�1N��޽4�j1r!S�@v�=���L��.�͞��0����Z7��<ğ��A��~,�Q~{-�K��ݞ_d�* ��B�C*�V��Z�����i}�L���z8�ݘ�\mh�kp��o��-0H"�P���Tm��|!�<%\"E����Ɠ>�cۻa^�/�H�@��LT~�Ud�Au?��=e0�%��f�I�{_���P�����t½<��.H��4o$C����YT�%U�;���+(�`-��4�� ���Ԇ���/w����_!�O�]���te�= �!wր�[�{}����n�ҏ��CpIJ+��K%��!Mw܏�3��U������Ʊ�0;1%r�Kl�Q݃�%�����_\����\�3��"����he��*iB��Z���S+�:	9�"���K��������|V����Yp��Gɖ�zi�&�p7(�y�}�����Z�Ĳ{Ӟ�����VZGƜC���޺�3�Ң ���Y�]ig�g'{��"5;�Y��4��?�W�1S}I.*��5������>=%��&;q25r���*�a���ٍi����P���`�p.
Z��;Ls��mӉB���H)+��4�e���~<ݢ�.��w|�s�cc�W�x-@d[�Je�8��P�[�B����%/+�p��bLq��UE 1K� zD�k�p�F1�qs����7؞�t���~
٣n67��D������d�i#�9��4r~� ��/��{�ty��v�	_ld����oao~
�2�gm%M���x��Q����'e�8�4����?0���d�=�ok	/ !�$�=���t��t=�Լ��=�Ah?rU$8@��IN	?δ��_�+?'�[�u��p�a�[%W�s)�� �t��;�g�A]0H��I��1L��	B��Y��pSXǠn����V�-�D����*O�+�ĺ�$[��3�S������Vs�U�_��p�����?� 5s =%vs��F�c�=�eO)��Ϭ�4M���7D�$dÇI��V!�l��5wu�L7��B~�?9��٭�](<�~����\Gx]~W��
�4-ʗL8}L?]���J�}�ҫ�ʖ�� Z�r����U4h���vy�p��ҰX������i/��-���<ʽ&ieYI�$��R�z5��E��cq�u�|�N�/�?̝�i��xW�C�@�,�vS=y�<�'�Q�7�{�j!Z�
����Y�R?����h�s���N�u���;��7�O��I�t
�T��:��IlMe��5�zF{~ ��GQCf��x����2���Kx[���%ft�����P*�P?JBM~#��*�C���¡�:�"8�p�j}�#�v�6�0�{�>>8Г�D8w;m�n��~w����_�n%C��糗	@�!�b��YO\b��Q�%���"~Z��g����Ve� ��^qn��Yp�W���9���X���@�]����=o�?�k��?V���ENx�'��P�c����柑�$��w��N���9XR�(����R��K��d��L��k-�}5�3;�%b�N�'��a�Ь*��`�sp/�����U���2�&�3\���r��*��aK�krָ�W�t����K��t�i�VS��k�Aq����;�Γ�`^\���<�f`�򜊎�a��mY61�Ѣ�}���j���ON_�R�#������íx˞0��V��|�4<��m	��d�~NSB(��1��u.����-����S��*β�@�
�b\�(����(��u������Q���7#s�"�	���M�໙5?��_Sś�Q���C�mq�g
�]+�0k?-��,�j_�	r����?��&".�g�q[���U�|��J:|_6�F��tbcp�z�=����[Ȗ������y�鶶���irC5�H���
��{0�c�Q��T��O8��ukx�m@cd�O1��%˓8��
Z*n�%b���1�CjS99�ef���M�_=R�r�ӵՖ��q7�L^IET�B�,����f$�.�G�s0�b�$�*[��$����f�/�SY?|���:�9'xv��@C��T��@��s*��	��D0@A\�l�U���ڊƸ�_�mϗ��]j�"�Cɪ�曤2l�@�4�+�R���[�����]����A��4Ir���Fǯ@��H��!���I��?a5=�X`�9�J�QK�nHmc��H�ۗC����[cg
�?;��9U�6X���xZ�v���i��ơEx=�Mm���n&�����-�,�s����E�T$��U+>�`�d��CP�Z��E����!�S"�}�l�8��LF�'8v6��n��3�p$�Y�Z��j��F��HO-33���ؤ5e�����p ���|���~�g�E�S+^(Z��qE��꽣O�,9���e^�[J�3��!��Rb&�����>�o�pO����#�M/�Y�{���9�]��+s�y��r#����ť됅���#A}���Dg�X"��7P�R�t/r�7��0]��
�XO��<��o�TPI���	�����m$����s�ht7���X�'F�Szrl�4"�Y3	�mQ�����,�ʿ��7��BW���~�c�[�)!��ū���`j�I����%�^��O]���b�M�3>r '6�%�O:P�� ��p�$�aW��Y0~U�Fr�����lfI�7ioӌ�fz2-��7����q��TF9�*�_��{�Y��w�-r^��
ڽ������չfP]�cQ��jBRҡɝ����#�q�,��`�S	��~�M�v���#G�gk�& ٬W&�x��G��ViXl��1o���kű����<�2��cZ�:o�9���Zߋ��(+f_�gx�2���m�Gu?É�=��- �W��۝p�
bX�B���C�hr��7�ui�#X���v!Ｖ6�vA}`��� \���P�\��79*���9!���ڥ1w��lW�h�f����c5Z�{���ɿ��t����P���=e�w����' ����f�m0���r����:�t�i�|+ŗ�+i�N��*>[��H?P��=>������9$X(����OV�:d��9�R0VK�[nB��qu���pq~HD"��Ω}���0��@����y26�-#�C�<	,uf�꘿�o�1+ `��u?��z�	�ۄ��F�56ڮ�7M�W{��	w�885B�N����*.8�i��v��EG�@3���k�͈CFf��"����֘��-2hҒޑn�)$�O��3=�Q�߯�"�j��>�P���O��#�H6��,i3��������<���<��!�����[l��D/@�YS�$���%�Wt���`��g��[tB�83φ�x��s��]��i� 5z�2�}��V���-]0C@��=V�Q/��!�>O�1�l��bo���`QƊ��#!�Ȭ�թ0>��1�ѐ�q�R��ϰ���0���<���3��=�>����d�XlxVHYEB    fa00     910�HB��1�f4�=yiu�1
3�cl^M�P�vc+s��Jl��i��9�תLL%e��?�֘e6 � ��}���+]��|(���m!�u(Mg���7엀�����Ǩ�6u��F~)������u���umں�����vF3��)�0a��=e�*��5�]{��5M����K7#�o�-����ڷ���Sd86�K���#��O+7�~�+n�5h�V9��a�|��k�u���N�l�3ӪTIs�hE�f���B��@�N@�Ee*z��/�L2#��)d�9L�cCov\P����*W��s�K�>+��U�b��-�C:=���!׮![Cc�_��$�vF�u������\(Xk_!HN �}e��w;��H}���h����Us6 K�u����Ǭ�bp	'��Ӻw���9�d��l�9B�]	�G�;�V*�� �eC������m��T~�C
ԫ����D=��h�EJ���~�<�����[u)q�e����=�P��>�����Z�F�p�c9��J[�]��U�ҲBxF�H�%
N�)e u���o2�Ov�`�_b��P�����O�� ��@U�g� �]�eƇ<D�b܅)g�|"�v\�j�m���l&���Z�O�È����p�I��߀"�Xl�l�+��j�kz�k��>�ˎ%��4�؇Q墨�kp���3�X����@dh.�`��U�����8w#�X��Ю�(�<�Ƥ2o�׿Z�p�O��4�"�y5��yy��8�������_��>:ʐ��q��@+�J*�_{�%F8�ϳ �z���C����Za�*���i>��W��$�8���u�����k�kk%�7���I3���nضe�Y�rru�/�m��Ee��?�6oM�������Zo0BSp3�ui���ޞ�r��{�z���:��bLq���k����\�2��{D�@��%V�y5$*���2� �6�A�U�*��ݫe��pM�h�(�"jW��~�F���a� ��7�)�̂$W�D�����Y�)��<ΟV��q5Ns&W@����S�未�>���<w��iV[sP�����D֬.V�~�T y6��XX��żzh|Ѹ�<`@^x�NS�j� N Ћ�a06gdHS��X�7���f���Hؽu���0��z?�����Oe�0(*�����Jf����᝞\�(X�e�.�9��?��z=���#�b�]�Ob$�V�ch�M�ϔbү���h�D��6��/�q�^AM9b��`oL턚�����a��8"��#��e-0��+7@�'�Ct�2�ygփ_����#	 ��U<��"6{i,d|��OcK�
����,�� ����Qm7/=A��a|��XpliƯh0�[�4')4td�b_=et�z�F'�1�_����Y�EK�lTگ�#�����}WMm�<~�� C��>P����e����jd݌ii�P��ljuo�6E�`� ��OV��V�W��m�-(4R������g�'��Kf�p���g�N�tnfA���D���A��Я��)� �i�K����E�mw��%��!���ߚY<`��?���/�#���n�2���� qݵA��n�Ө\��,2Y�Э���,�a�hS0�<.�̵NT7!�<�pT��)0���ۘ�[&�:
�Y#��
�� uT~mv+&%C<�X�#���u��0������s�u��#̔h|�A��z����ٜJ��_[)��������Ȟ!2)g�p=u�_U�l�O�p�C{U�篑��Xs�:�K��L.�ƥ �?����O?5YGP
���C	��҂D�b�1S+��i5��Ί\�/F�R�lc/�d�I@�rim������)��|(=��� u��tmM<�/ni��%��4��bith<lGu�s|�j�	��=v1���ܳ�M��d�J7�n(���?۝UAU[�n�Ek�e}*��+>P��J��3��plRM�l))�
�t�}�UXx�3u�!�bi�Z�Q/�r�ـ��J�R;������_$�%�0#�uTV�w�E�4u�8�Jν/Q�2jz3�Z�>fǶ�����R��t^���������`�A�;XC}�I<�[��"���V��!P[��1�p6�SaEn(��k=����e�#����`�
���SZ���:�z<��e��&� ̦���וK5J�0�,<q|�7�q�$��*g��jr�\)Ib�;�H<��o�`|�Y|��}ԼH ��σL�2ht�j���&�<���ѥ�k� ���5��jXlxVHYEB    fa00     fb00Rsxʀ�s��`������O�z��7���r�Y�!�j���J+6�`��k����#�ҫ��Ҧ���+������/%k9g�N�s���ۣ�ф��}�ův[��&g� r�JR�p������aM���u1Ǫ���91��A�����6��}l4Vld-���ɎK�p�B���Jb/9�}�Cn}k�X�
{�G��J��S9�,�?l�L*�@̯p�$Ͱ�hQ�B�6@���<�U�'gۖ`aY�G��w�!�pP�\T��*h�( ���%uÇ��0r��|�-bؓ����-�$`PP�K�4��O_��M/�10��-��+�y���T5C"��aQ��U�[�>@)wVdvq�s���,����{˕��i:��˦��1��}s���#�u�J\��8��૨��OY;���s����w.��a�5��ŷR8+K�����E'w�N5�j5	�P_o�����%�C�|a(�q��=��N����f�#���¿:��u���d��w�u�_��wňu*�sS����y���<�9?<;>�ڰ��,�ĚQsl��z<3%y�:��)+o�H��rfr��<��c/}����w�ᄪ��Yl.2DրE�g~,��qx5��;@�	�c�� s�?�l�
�&I����#�8!um*�i�}�_� �?���oyK�$a'
�K�� >Hp�o�H/b��-%�7L�럭$a��t��#kq�@�D�w�j�����)�~g��4���� ��	ԘJ�Q��h}��<��J��b������T�=�{�[�2..��u�[.K�g�U;�-�P����pE|�꺲���PZYe>adK�eU�'�L�5d�LƵ�#���6Qy[0�cE]��I��U*C��S�^ו^r(I�FT$�`�櫰E|�.�=a��bRӗ,���?,My$Rn�{�v#m�k,ʇ����v?X�GeZ�����oL��3R��t���C�)p���Ĉ����r���R�עe�C䫖\�[�׹�]
��ݺ��)9�eOz\ꡑ�dq�o�^�Z@ɭ�S���j߲O�9����s����>d#nj�jo\�^I�R�0T'䕒�M���DD�b���gh�lxt-�ƣ�E�>�̌��e;(8��������`�+8_���#�#o�5��B�i��ȁ}�B��E`�\3���e �}!�dZgi��jK�����0/4�B��
 �"��
}~wY�(;Y3�/�˂Y|>�6���Y�T�O���_~����3Hr��<5U���uRR^?oO4�)�YT�ȇol|�5i�7/J7����@�zH��Z�jvϨfh{,��u���'End�A�ŕ��}��]�#�|�u�cd�,m�4 �YW8oh�a��g�n>�Ȗ��yn6���?��M��q��-_��©z�E�w\�+���rJ`|D�����H�l�;6�F�CD�2���c�#�-x��3�:L��@�o����m�A����؞�O���s;�챻�=�nVJ��đeZ��vɸ#�"�_[<� 
9������Cǐ�����	/���+!f7��{�ѷ�(9�5�X�'k���̖�"��i�6��s�ڂ]�PC�ܽ�BwRȌ@x��z=��lz@���:�;����ݣ��� ��͝��X�"� ��5�� ��a6�
�%ҺVu�Ƅ`4�K*χLw0��Y,��"}�lً�=��pÕ%�vi��%Dg���,�?"��Y9�F1z�9��*���TQZ��#7��W+�2��M�]�y�X��M�U)g�������/^s||'���/����_-L��k}T�������'�1�KǇ���Ɔ@MG /���{�{�v�Sz�:H.��ʾ&T|g�xY�0+���x4`LT�Gli�ս�"0�����G�P�wb�P9׀�3�]���?�h_���<�
.�jQ��ہBR��7�̱��H|Qf"zTj;w1���Y���������b��I�H�X��&x�T�,E��x�J1���!��T����r�+�^m+JA)������j��y�
cn�{�E�(�g�%Ą'6������֩G�&UnT�%C�2Y-ya�g�_���ڳ�f���׿Q;�6��9b�t�k6��GQ�~��5K䒗��	�w�Ξ��6Y��{�"��E�Àx��k=�0r%�ߜ����j:��їU&����QD|:	*��!Oڮ���|lˤ0�?��0Q I%��a�=��#f�DmxjI��=���\�h�,͋�ӗ��B�S��+���R�Ѐ:���$ԝ�|d5�6�H�K�4�LJ��ǻ�[�lKJ+��#&()#\�18���z�Z���45O��ߪ��ɂȨ�O�|CAz�c�N��nc����U$�i��&�wmU�^�������(�!2�9t
_�����aA䍫0���!�η�@ ����nĞ`s����У33TL�g�qJ��ÍڳGf����Սlh�I��*�E�<���p�	껃���vE��Y�vܷ�r=�YoG�y����(ձk����aʡ[��P��_�unw�:������=�4�EH �U�z������O�����ա�3��?��c� �>�{���?D�-�t���s��Ō��A��8�.��xs���]|)�=�_�[������%�X���{�S�9���y_� |��^��H9�1�{xh3�L8�9D�6X�Y2R�?y`"�"�b�!B��%�� ���W�Mo%�ؠ��Ћi��:�	��vQ�K�� ��k~�9�r~^f��$�"�!.R���Ҩ
����Gt�:b9��s�=��t	���|�$s�-�������:�:Â�d����4�W��@��{H�`q�Č�	&6�6݀LP�s�K�h#iQ0T�-9��0|t�+���٠Y�x��~�6b��P#t�T)�ʱ?o�C�H����G"j�SJv���C��(o�畭��16*����4^V��X�y��.έ���vHa�|�z�� ��;����L�{Zm��ߘ\�`��e�����M-������1+���,�2�ץY������a�V��J��Y���z�5V6�k�M,�Gc���	UQ/v�~ ��ľҽ �Y��2�8XMG��Pm�x�Lf�S��9���]���A�����"T�$�/�P��X��i��A�X��ic��2��� �
��L娍k�P�!2��(}�I9�Z�ѹ,�6]	��5�-�J��xGa��x�@4�vS�ݩ��]�ǤqTM�s^0�����L�9QN��Wf�S�g�_�T��}�B�< �+�0}a�LƐ�+��=��"�MBTn��yj�n��ֳ��g����4�[���������;�ߚ�UO�>�C��up�����`*��&��ꊔ ��i�ɨ�U�b��A������B���͙�
C���E	��/^<�<�c�++�d�16[x�`7D�8�Gy��-ӧs[ㅳ�U!-�v1ث�s���윔b�d�t	:R����E5�������hI����	�;^��ۚV�_v�F�6�4���Ki�	:���V�Kڲ��V�~51Ez�C�CV1��}�A?i*�=�߉U֪���e�3
N�M-E5�c �`ρK���dH3��@��qZ����h
���7&��#��1$`7���K��-�����n
�z����A������7�V��p�d���� ��1�'Ŷ[�8�j�86�����ׯrv�px ̮R\�ǃfm�J~�g��cZ�$��liv�+\/�5*�{�@x}�{�?:8V�JW$�$1�CZޝ��܀�eg�A�������s`X^�k��ƾ��3��΅oM�1(p���c�AS����{�pcY����Fذ��U���}��Y�:��=���hU�uܩ����� Tߙ�[�@�T�}��H"��\�u���H��F�V�3�/A�K�z��4h�_���$fx���Q��XlxVHYEB    ea85     fb0?{o%�D��ƿ��.+-��um��q:�]��!h�@D��xF�#{��d�uM&��)~��yֲ��D�
��P�n됈��-\G>�{�'�)�Q�sȢ	�,l*U�;�TW*ј�.Y���J�K�E�Q@�}��b/�fSЧ��l$��Q���WK���򘲩 P�Dk��o�Ps��n{hϟ����y�mʜ ��0�$K|����K�N�L�`H^9_$3e�;ٴTp���'i��� ���&LQ�ƻ���X�"�z=5�WA�%&�skI�g��=�9�HI T:�	!hQ�����{��9�'�ڈP���F��E����h�+�vt��S��b$�����ʎc޳I�
�5<�2��	�m���N�ᤊx�7���#���o�Z.�pe~dj�7'����|�Ek��*�=�Y���]ԿH�J�aр4P�:w��v�����"�"�^�5�],�Ԝ���S��W�� ?��"�~�Fy�j��sA	�4�wH{��F.�E�����U���8y唩Ά��Y�2_�g�T�g'h;�*�V�A��jCGZ_��~D�͸��mç��f�xmU'K�f�+]簖�1�	$:##���vB�uAV��c��X\wy(���{i���7e��}�<9�WT��.3����zN�9�׃��%f�(~T-�BPs����Qq�j��i��� ��?{����˰ۄ�z=�p�\�� ���M��	���Խ��<��q=��
)c�-kTh��f[��?p��=vJ �^�m�=��I�x���O���-������/��Or���U�;"�c�BT���xW�{��-%����w�o=SYa^��4��ۧz��:����i��Xz�_Q���΢Lx8Z�C�q}��"5�U����5�p�M���G'/�2[�eLe��
>�	S1�.J��L������Ó�6���5����-VB�BC��0C<��E(5Ȫ���^2����T�{֩�˴e3d��5}�+�oJ���]��X�ΒԵ�i�u�3<Һ1z"Y��c8}�g��Y��Z���)��QI?�f�͞�JOz�ҵ���j+�u��ef��P�$�
&����\��{&�Ŕ���E=K�#��i��A�8o� 0f���e�R��jv������.����.��	l�	F�=G9h-W��j��VNjl݋/�c8T�[۪e���go�/�X��C��O�A�ｻԧໍ��UJQ�v�]������g��m�EK��Ժ�:HD�uKi�0�6[F��)9�W��0�|�S�&�&�d������@}c��YC��?�Y�^ʈBja��:��[y<�N"F/��)U�͞�+m�Hu�QV�Q��BDA�yL�����e��'Y'��pf��rA���w���iY�!-��iȞ�j9~T"�۷@n���sek�}�A��l_y�z���T*��j.�!Ż�E���A=�k,~��wn~�Y��� ˔!M��g���7��")��7{�"1
������&��Dx�=t��������(O��2A-T�AyU9���n��
���M�����ϗ� W鳳�7�T��:��.�� ����C'N"�{�Co����T�O�^���C/g@`u�*�3���Y��$p
�6�y���P�wh)�ȓ�G�[Lgp��ð�3/�:k%~��� �Ќk�7H��V6Pg�
o�&>�z@٥6�@�����N)/?����A� �e�]��������r!���#5	!����h9/�"a�D�c�g�V��Q�d�p[]a����Bё�t��S8��F2M���X�$+��TYI�֙�h�;��~�J���m��ݭQ:h�L�X�M��
-k����B��q��z�h��k��cE��1�GVU�O���zS<i����ޑ��hD�D��F{/9ݼ�X�=4�M5�I�Wf�gy65Rf?�Z��<E+��^��78@=�lHn@��nG��1B1*ܽML�����a,M�K
�%��m5R�-���U��Ѫ��7���H���*�����V+c:��ה6%JrS���T�\���Q�,?�R=��
�.%!���~GLQ��I��_|�l0���$�i�z>�>z�1�9��n�y�	��6�Q��S?Q���;�+oKf�Ige[`6���L<*�R#&0d��%�n�KŠA:ٯ�u�F�7���=��s�\���o���I-U���	3##��.��?E�^?�<^PM��	��� /њ���`��H��d1�w�Y�`��_��_�Y�r4)j�^����p?"��R���vY%C!�$�T��%�5v��Ӂ0Ԍo {'�ݽ5��>�������c'�#u����b�4�7�����xm/I	���<����/��#�w������Y9o�q�ZyK�	�:Y֊|A^�v�"����q���uY�6�Q����;��%�D�cv�$/�5Y!b!�$�rk�uj#o6AE�f)}KG�}����lS|�ʘi)��i�y,���h�L�e�Y��#V�����)`=��4��o<O�˧Vh�Z�^� ���)�q�d���=�����^��q#���^��%֩��\���cV�8�U=���4��ܲ 5i���@CӐC#�۠�7�$pM���T��{���TWۛ7�0�{���}/&:�)��phA��+�8M��DX���q�=閏�g��L*3 Q"�S��-d�"�j M`�r��6P?����x����+�;�V�=p����N'���̤K����n&�c�D9qwiyA�<�}���	��I�h�8�H����M�X>������oOE�{`�����=�Y���'�ZJGI[!�)�kM$�{O���k����u�;ښ���C�HFV������G#(|'c�s{Édm�5Jkj�y	�7b�dB��M%��r�i��)�#�������bj��p�����i�q���L����q�-�.%Ԍ]�$��b��~C&�=�>��f�Ҽ®�c�!��(@�}�r[�ZU��0�� ��	��zf��C��I���
��|��β��w��~�V0�4��'�q#���9E!�=zJQK�J>ރPKtO���]�t|قmI�d-@`R2^OգY�n���*�B,��Q���	�-����.�/Z.���)*�l���|�!@�$���(]�����~e�'�v���nBR��t�W�`4�s:��8=ζ^�O"�E���4�H����a������"�B�{4���k�����2 e�Ͼ0�r�Q����D���jO�����cc��[����M�����r��evF�IZ���؎�ڇő�������V�(��Hvt�k.MU��SB%�,��#���ī�u)*��0KM»S�5�y��������\�`z\�]�>AF�)HfT�2��*GW���EO�]�,\�F����tA�n�*���y�\&lsW].��c���d睖���A��S�k3��:M�_m���T��N�E��^O��p צ1p@��Q��䤡�x���Ky��rf��k
�b/�JLg�G�LP�;W�^|d��=oћ� 8O��?X� ]���!>1:��*C��4֚��8���bY~��z�~p�	�^�g�c�q0z4��n��<]$�)FR�x"�k��^Ӿ�x�u3���+I��٘ࡵO�h/~6n���J�%�v;R8�ޒ9�eh��1��&��M	K���U���G7�˹��M�)�`�6�fz�j��yɰk�����c��w"qvR�q^��U�u�d�j�ԑ�g)�|q6bU���Wϖf@�!�k�ӭ� �H(��+���_��u{��w��������T��͢���R1t��xE������i�+�4�j�"�#�����	�����4�n\�����l��h�Ֆ&�0��b�a�ێ*�2�^d�$[挃�{k��P���:�bZ7`��z�