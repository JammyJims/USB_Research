XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!>*��>t׶�KL��$V���э�u�,Ar�|ʜ#z�!A� 6#�@DG0����'B"��n	2/XZ+�o�t��2�i�r2�Ew
n��)}�����#�ن�;�V)����k|V�p��a8�)m�ʂ��纚ԅ+Ĉ5	~dm�d����[���O���T�lGt}W���2�#q�:������=�T�E��Ź?1����Aˍ~���0��:�q��*Lg�S/�O}�z����Rב�����LKm�	f�	��Ē��S1WǉNp�����nUqXdu9ڽ�����xA'��HJ�'�M�� +�mg�5��\��>�Qm�ndQ~] �-�[�~�T������ˋz���9ů��-Cdrҿ7eC>��4$\��g�$K�|eC"
`��c���@��~u��1� �`Cn�5Q�B�N��\o��]��<��y��ھ3b��$*XF�8���yՃb<��8@w=K�a��	��9p��Af�F�m��o�8�`��r������7j"1A���D�̔T J�B��9y֖!�,����{��2���&��Ë	������JW8�l�z��x�.�J	����S��S�}�n�[N1�~[��q��;�.�p�R2����5U�2�����#�����q��j���wxE�2^�<SK��n�Mc`�m��l�u	
	��9hĞy���ݓ�ŚV������U]oT�aa����ֵ�[�ȥ� �+���}a��E>|�qMSXlxVHYEB    192c     850������eV��
��M�ZX�� cNk?�61x�r@��جS�
��yq������6�e�#���H/0OJ,�@-I�*lE�ui��S��'@"��5 ������-��'Y�p>�c�)���\�;İ=�v��r����BE)m��`�[;H2A�S|�|�b�
(�.<��cN�qoP������k5ڇ<�nPe�	�ޯ>L��"q����.u>�_3ʩEz;�|N����/�@�j�%�W�y=��X����'��pk��t����/���0��߹w����,.�/�o#�@~�k���i��֓��ޯ���H��o���_��bld�[�f����H�v^y�Ż5J�s�*P?"�.؆�)m�63��h�r�lf9Ү�N�����l��p��C*�q5��2#�����YuȂ-�����옇#m����MN���P��f&r'�	�����ά��`����e�[�H��M���>%!"_<��r)�h�O�]�<��r:��~ķ�YA�x��|\������K"�im�vq!�VlDz��G8M�̻NG�u�!r`yo�[ѷ9"w�ݗ��A���!�8�65�#]�#��v�p�P_ᇜ���Z���ojZR������s��k���Xe}%���k��BSE��H��$v)�2���佭�E0t;l�G�.��w�6vʚ5���F��) `���Q��3�n�Y�0���f���=G��a�K�~�@�5.tbtBa�N^.��lW!�;�a����l�w�I�dq��tJh��\jy�Y�\��|j�N��=ut���B:���q��"�Y��!Й����3|�.�Տ����a�z]��4o�5������e���Ck�R\����(���
xS�}T���-�
��X�2��}z�>M(x**K>�;� 頓{t���熂��_Ak-E+����'
y||J��kN^ˊ�p�3�b��+l�b�Z/:���ŏP=�&�6�Lћ���:>�fb�^��2q/�t�Ee��Y�VJG��u��� � �V.+�2�����i�� ��C�I���G�XNa�%���]�]�������nq�t���j��J2�6ę��Y�FP���h�ݥS$J�J�f�r_��P�3<pSښwPTkᙲO)�b+$恽b�5d����ɚ�Ż6&ڬ�)����c�����=����j�r�ӳ&����l/�W�h��V�932@���� iФ��l���7s^�j�"�vq3M����;��������s`�d��!���98�:^>�uM-�g�t�+������H���-ۂ��Hv�ƹ��̚;nm���]!�H���;F���]��t�kX�UȺn��ϯ�J���5�I�ړ��e�)��i�2u��/�I�F�,׵y⾒�ˇHg��/j�?S�aKZ>�L?�N���}�O/�R^&)��yw6���˾�[�e�'4s�݄ҒWa���l������9^��4�d�_�G1%�P:K~S�.�R<89�;)����)K�X6���UG<U����T�t��:�rZO��ݶ�0ب���r��3�2��4��G�Zm��9VN���œH_אx���]kt��ǐ����;X��׈l�g���p/����I�#xܱ��ŋ�X~0�OQ+"�cȻ�\w��Tw��<�"��^�!�=)mkN�o�Ac��)/��pn�ٶ�W�)�$)�!yb4� ˡ5����)�:vs�̈o�R&L��/��tmI��'D~�Q�T �9<�j՛t�;N�&JaS���1=�:�1��{d}A�>��g�_�aO0�k�1m��[�j��~�Ŝ�wc2ͬ}�e�[�_���;��w��M*ض)���
��SǢn�h虞\���{�%m4�&Ω��O%��o�(��"<ʋ%t�~�J�Sg�8T�/���㪷��-��,D��[��\p�uo���C	�f޻!̤ljR��;���'�_!�vE��߮�Qq�	�rvx�w��A�.Yڭ�͜���Q��ޝ�w���n�[��(ich�ƪ�c�X��M�5���a���?Q��jDīCK�(�L�,��V�Ҩo��:�\pڊ��