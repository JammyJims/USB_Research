XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���cM�;���M�[eTN0�:�S����E�Q�Iy�	�
�}ٹ�pYЦ?8����*+.5>IC��7�
n��u�����(��R�&�T<7�i�z�m[ 	���o�mgZ7�`�񆌂l9��9��4��9m��΢f$�n)��B���,���.p�U�eЪo�6h��Q**�㧋����#=��0�i>��\�d)YZ{;���Y��&=��m���׎�ސՖ�.�;M㙘�D=&�߻�KKK� ��\�«-������0��뵭��q��H�y�&�I���]	�#�
;�&�}0+����o
�l+��C�jrdS�O��
���5@j�ai05�e��C�Z�pxV���U~�����U��?�59��7�7��v��lB��@u9�`��k�������l����HE��m��G?WQb�f{@h{Z5|�r�l^���ˍ����L��1���J�d��>�����-[,�%n���H �b�������R9����J>֮Cn9�ٰ"�J$�g�=0��K_���ߏ:�X��S3SN�7mgᬫVU����:f@�q��!M�χXQ���~H짒�7Ef⡖d#����d����ӉH���"R_U
�	�{.D�w��0E��-hxf�<�W\���)��3Rɟ4uB��ŉ���F�����(�����P���E9�Y`B\� ��\��@�9��פ;��B{d�i��/�":��>m�
��R�1���J�4�h���=*K�XlxVHYEB    36f5     e20���5)��w�LQ�7�vb��v5��J2��i�ح&Ү�ʐ�VЂS4s�e�9ΩKx�Nj�9[+W����`��G<�3�#�`PlQ���R�1���uTcJb�C�=p�v+���P��w�mwH�7MiR	^�mQ�e88E��
�ȇ��D�?QZ�W�Ѿ
����Wۯf.�/q�䄎taaT[|��=8�qM���v�_j�z�ɻ\N��NR��MU������F���9�����(H�9�
�ʻ%�;����9:[��C��![�C���7Wr����-��ڤ7�dj@��=n~��ڷ��^M�O������(TB�w���#�4XP$���2"��\���>�� ��8̕x �Y�\	�]Щ���ˤ��sN���,am��gF8x],�(Ǚ��C�Lg�U�I{�Q�93��h�����D_��6�h�|W�E��V��b٘�|B]7ڨg̮�\>���pe<�\[�5ĔQ��[��?&!�|A̙�!T�o���������]��_i�Ǝtz�
���'R�픕�48���!s�I7/L�Y���O=��鹖�Z�QV�5�A����=ptvD/�ƈ!I�J؊�4��5��H�Iu��%�� fʪMj��	�0�}#������@��\�]��#]�b�c׉A�A�k�s�:�<!H+N]�ƚm��Gt��OH&�<j�����P�adr��w��Y��cǨ�������8,�	�֤y�6�a�M�S�U�u����B�Wlp�R�ƣ��:�?�lr���;�.�p[�\�U4� �$8g��j�c�b߰�E��J�G#E>��WH�֏˾�HX��e\�ޏF���%Z���Ԍ)N����]���}����\uɃ�xqd�
���	f��<��̅�ih��{��Mo��I1h9{��`�}��i����w��'�yFՊ��2�٦��K�8ʐ/�]P+��S�x+��a��l�H�G�
Kvk��OˉF_+�,��`_�%�QC��>�E��N37Χ(D�wEwb�޷��H���L B?"�yJ����L�Ћ�:3$�eC#�ˉ4������Rr��� �y�NI�+�p�*�=���A���m�Ѱ�������?1&3X #?�������wTX� v��Gx�Zl
�lyF>�}�	� b!B�8\�����Bh1�m���"k8n���J�a�_k���۞����y�w�����;���u_�7�O�h�H��z3Qq��>׸�$���Յ�_�M�>M ���L�� �vh�R-�f#H�z,_�a�����h�X���)q?a���E��#m��P��;��J���hɣV2��4
CF�7�8�iՆ��7T��V8�H�����	���e2�ǚ?K�1K�����x�ǈ���[s
1r�r��s�C�R�Txalh�8a��-���p����=�8Sˌ�|���:���SZQ '�7�@ %{��������Tr�շ��Zj�oE�J{OO��F��2v����.D��^y??J�X�6_b�$�q�����X���2��n<9Ǣ���IhJW+[�	��1�a3�\dM=8ߧ����PQ��)�k��>I�|��k ��D[���v��+̲۟*Od�D(�5h�d ��/6�ű"� -�]^��J�K�"%<� }�ӧ�Hc^�y�����@&:�q 8]<�)N��6G@��~QA�,3�����Z����f�ͼ`�V���=}�l�OiL+���Ͽ�S\��t���r�������X��
���		l�u����rz�V�O=��އ�K9�r�Z�m?lS���aK��݊���0��QJ~l�pu�z���w�Ѽd�8r�7�ԩ�[�'$
�F��;�[���8�]���ݝ2_����?K�oH�T)�<�{�ɖz.&B�cL#���L��m	\�+ؼxf�|X�D�{�L��/�kr�!����#�]�^���;%�F�0N�?��&�u%6�G����9&�����FV�e���x�9t�>|��K��oz��[��1;��Ӻc\��9y������5�A��D���0Z�_��߱��y趴�"�!�ܠ� gW����P�d�|s@���;�O�r�C�*zQ��!^Hva�2���9�x�E:HjW��j������#q�(|����q������.���
��t��2HL>��Ä��\W4J�	ȋT(�wn� /EN|�<�o������z
ò�8�xu�+�bj�\iB����J[*�O����B�����k�+��?���oK�<�-�}�I��aO�L<a��s*m��RyI��<��A�)�R۷�ЖtU�5�(g"kXľ옏w0���w� 4E ��uhͲ:#���XK�d�|i��Z��Q�ڙ�,�T&]G�� I�L���X ӗ���9���s༎�5K���o^mdYp��
4�ש�~��B�%���h���W'��h]��g�@=�Y�~��lΗ��#T+�i�젺���]l�-�ux	����NL�(��
�d�TA�V��բ�P�7��Ȉ����/����Az���R�¦T�s��5��%��NJj�4����JD���� -;~���r�O_G��%�[O�q\~�{�Ί��#���;�K')�{i*���Dt2Y1��ƕY�?��/"�^�&�t1o��D=�,���b$]0R�PD�K�����'o�9eJ3[g���O�:�MB�T
�|��z^ �$9�ʉn��9^��B2E7������@b�AgK�M�l^.&��J��s��m]ȯ�C���`ױ��/6�,L��Aj�G�7�K~1p,���8��]YC����]�����l��q���S�I���M�곩a������g�]�o��q��}p�E�`���-	a]s���ֆ�� ��	�%��c�)��_U�1�m�W��U�f�K�u������Q�/�+���Q:2xR��%\׫��hE~�K�܈�lu7��5�O�f'�3�~~[9��H�E��aΘ�& ��1�M]�S�Wpd�w�aal8$����
��ǉ��N��Gz�>]&Z�k��(��t����Ǹz�:��_ �vD�'���{O�'��on�k[�q�'�p�2����@E{�&_i�ef�N���ݐubR�N�4GA���RbI�5��ށ	J�l�����*�>[=:,'��J��3t����O����n�.I�3���On���>�W�^���^N�j��!I�$�x��{�)��Q�
�)��d-�^��E�I�/f��|��U�3��MI~�ڥG̹��=	L��:�Mȯ��*o�N�J<�)�����
����A�0����/%#�l,	@?�{�;����Z��EԚ��'�L�0����Cx��)ǒ�ފ{������R�겑����?�bc��(�7����Ǹe�fxCּ�2�P��#���b�v��~�0��k���$NYm���bq�ԇUЋ7a"PP�0t�><r��#ԏ�A"E#;9���'���n@MYZ�ց>�;\+'L�6��_m��o�NQ6����  �cD���*9��L�|�o�D