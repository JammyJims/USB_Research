XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~h��Jz״�\<?�9օ^�C��X�א�T����9D�S�KSݐ�� ���J�n��^N_��gh8l�2q�2>���)�"�C���*�}�aĚ�@!cY��O)�S�lxE�y�; >�V��$�8���;�Q#b��%��6�oդ�@J��_�&�����H�I�\d����9{
��g?�_���o~:�@�Osћ<�-Nf]�U/��5B��߅���@�J�{���@�┒SH��Hj����|�p�Yp�r΄��^[�
?8Uu���wǴc/l��f�X���o��M� U�����Sq�:�iY�ʟy���%��XO��dw���z�n�����%����{�EǇ�sR-����=y��O��k�H����e8��&~�K7�`d,89g�:jbÈy�H�*�y��{h(�'�	!h"�<���vO�Lk�+w�c�r��A�o��%�;��X>�4C =��8�gS#J�/7U'�<��U�3_��c�?\��S�'�U77�v�ˋ�\pe{ \e�f?fZ��ЋN����ƅ1\����ٱ2{m����-Y;�Ⅸ,�o�uէ��"��9A��Z~�k�V7ˤ�C2�e:��5�z\W �|�?���8�s����i:S�9��m�I%!�)�n�9���8������iHⅱ:��h@�sl���G�;��\��\�u!����mB��������Wu(�-ty�N�0T�|0j���`8Pn	�*D�Ԙl�n�ےx�}��-E�D��k)�8�~�XlxVHYEB    4324    1010���]����l��2��s ���C)v�X�LJOS �U�]�4���3>?
7P| ��!�ޤ�c���f�r�aE�*�U��>�"��IpGxK��a�+����������⣫�\��GtQv1�p\q�H��M@�Wm�������=�S�ox��̣B�����$���(flL�b��v =t�v�_=�Q\�a�v�)l�'��<,Q�Y��)+8���ǭ�����6F��K�I���N�r�E2rU
 cq��Z�b^���:����I��1��k!�?s�H�kɢ5R���ծ�Fu#�6�[Q���_@w�˗��,�]�;P��ܾE�)�i!�[���q{���6�Z*��d�O���T�ۺ1�KC��O�p�o�q�o�%�=������G�%��`���RrV{ۜ\���c�CŞ����jeC�Т�;��Y-  GnZԸ���|�d>��`��'>^���3Ʃ�([e�"�ߗǭ�ܾ�*?��Q95���h������G=~�1RYdf���r�ѫ�Zl-�ݛC*�g`ɛ��)U�R�f4��Q�T��FRƜ��)L��%Oaa�e@4��Y�|(�O��ȱ<��c�LkM}d5M[<���u����
��}>�N�l:x%%��`�w���Lq �: fe*�4:#���H��0�rF�r}����B��K�2��Z�qHS�."��x�p|A�M��� Zf>W۬���
��;�@��G��E���T	��vq��D3H@�i�o���hNh��`k�Q�	��@���^@6�B���؉�M�[.�y\S^�jo@Y��ӑa�}���޼lBVFbtS�!�衭&��p����M�� �]�[�F��>2Uh�up L��/V��E7:�=����ԟ��-h�n�� �'Q]y�ςic��Ϋ3H�B��,�K���m�.��q�g�ƐBLo����0]C���S��o�I՝�9~\��LY�u(1����.�#+t�2�_�"K�4d�1��W�Űuˉ���]1LC�_�쟼�x	��l�չ�He��n�{���ΑY�sp?8~���=3.�&��(jvpv�F���\� �z ƻ�|�����Z��İ�!1fr��^�`BE�@���~��GZ��"?��M�݆��M���/t���R��~eY^�M�8�-EAs�G�äK/C
�s���p�q�/���=���y�y׳�ujEV�ҩ+2��=6�� 	5����l�Wo��KQ�U�.�[�K��'�D˃�g�<4JV��n�%ʒ@>�lV>X��A�Mm�%G]����-�0 ��P���o��W�zY��<�4�>$��;  pk�sY�Ob:�6������_�6Л��)P0��Oo���=�`��9�9 �~�f�� ؏nʗcz�"Š�A��,F��W�8t�R��^��/��yiv.�Ѡ�,ݫ(�L��yQS�s@��c���t
��#o���0��E�3��C�]�Fe�ɢ.�tL���^�]1���$���r �7��~���A2"h6aX9�[��f�N���ӭ9 ���/����?��`�A��~p*�$�	����w^o�'�cG}(����W�u�*��~�Gf3%Q�Ͱt�D<��ƹ�DZ��&�����#��&)zS�x�F�5�9 ���n|�=�r��Y&
0e�a���(�T�| ��Y{`�|5��u=�`@:}�P{�Z^՝i��~�]�-�??ޤ�n4�fX��+�����Ǥ�6���:+��>�����ʹ� \�Gr�ñ��<k����)�4��e/�	}�_D�Ӗ5e5������}���1qz�Ӝ����PE;e4[0]U ߶"�a�������FY��[��\���9/���<��U��b�t��&����d�ʀ	s�_�i���<��-8xS�E���9�;�����t�g�9h0̅�W�X4��)��F����єcyatK��#u�E�=EԟK�PY�7.C�Gy��@���!Q�bd�C;�����^'I�����>y35{a<><;r�G�D
d,���\�c��|���b� ��
ۺ}�C�T��p��?P�=򬸱���
��!�N�"���k�qj�Q]�~T�	�78V�l�A+�?�p��g�L"�$!$�ֲ poCZn�x��j�4(tZ�5[60'�xǆ�ǺGN���k{�A�Z�N�ԥ���s��.D��&�.����H���](����@[}dQ7Ǆ�{����c�q?��2M_��o��`󙩬v��g�8��@q�S���捗�\�t���B�PI7�e��k��~��h��A]8���G��`O��(z�h�.iq��8XT���CSa�Y��xB$�?���f!Z���W�+<Z��<���$��x��^Xl����>h���\#iO�i������.�<ުSւ�nY�c�坂��w;%�7����s�%:3U����p"��'�����wa�%0�|W:8W}�)�N|�>�hJ��f G�c\E�&�W�r�Z=:���*o�8DB���AuϸC� npMj��1����2�z���^�JJ����iFW�&��c[u��~��s�
�	j{mݽ�(��^.�9>CTܥ]�I��8���+�q�*�\�r>=  }<���!���d��d1TE�Yx�ey�u�!"�U!�GŧyF1��5k�{R��1���ܾ!�Z�9��r�8\���/�-xxQpk�O1A�c�h!C�S+� x���Y���3r�=tR+��|G*��R��5���.�Ģ����X,+�"h�])H$�)O8�g�fl�3!���z#�a�"
�V���:F�S�2��/�S�	��"�cC�
���s)Vu�:bw�įB'�r�D��A�`)��Y{�^���1]��vW����3��1/1��؀E�T��E�I����.�x��aj�}����B�CEZ���Y��!���:�Q����U�������m�_Mzg69�"���W-O�C�ed��W<�����7'������Ƀ�-�1L,����)�f�h�Z�p(2�A�J7�Fk�#����-���W�n��Q@U�P�4��mmG�EǼ��Ļ�S�`罃,-�p)^+%�ĸ��$�9p�X�v/�8	dƋ�[/HsM(D����*�6�?9����6��2N�Ba�f�B��S�kHc�RI.XO��_��ۋ����5��*d�Ju4��d�L�j;����5�ibS�}h�����a�w7k��ø����ZL) K�����wk4CrX�(i�Z���]�a"�>qѻ�)`<�ők�8��,>�G��[��X��O�+�z
)�2����[���2��s�ήՀ�ޕv��mQR��M��@=�O:�+�U5��v�}d�(Gވ+��V�E�y�k�Ð�: i	���Q������4�$Z	���?�ˌ��܀����҇���>��b�ʻ��gPB�X��T�D�fIU�k��d<la����~Y�:c��%نq����9k��}&qe�Fjd5	9$}�
o�K�P��-��ҟ��,I�����z��r"��X�3�S��]��b���7B�l	�Kvy�,�K�x-*-�,W'{��N`�Z�����'J��䇞]��V���c[�6���뽿����܆�,��bI�P�s�{�}�f쫛���ay��ק:���L9�sy1�w�(�k�|���La���#�rb`)�<-����(�e�Fm�y�����9Y�G�[�$h4�v~?��B(SQ�|�Y���o{x��{��.T9q�����>eM<����;��?|��Q��6,��p�UDiʤ�Hs��%;���4[{Q\a�]�q��%�n��Gr�UN:�l��JC��U7�� �w��)��ݾ��*��O����g�jG6*Zx�)�Fc��T@����;|\�A�{��sU�����:� ,�N<�!�1�3��}�lXڢwD�J=cۚ+E7�![�4�/D�g����;�����+D�jV��ީ\�#w6M�F��
�������zD� �p�Z��0؄g�߰���[�4.������"�s՗����}�5��>�% Uj8�ޟF��Ff=L