XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���k��n1�{��qY���l���$vZ�Gl�k��	�e5t�����`��O�6\d'�#/���k�_�|u0�7qvd��B������? ���7~֡O0P v4��i\A[��ԉ��m��l�~��leN�	x(1��%���	�D�Oy����hʒԘ3�5�[8��Bb9���C:���:A+���\c���6��H(�Ÿ��r@،�c����.&]��� �}8�*74;�1g��'s7�!����<��5��$�A��������'�$�� �g��!u�X�
��we�(Q�w����CY���}�>wv4=lNi�n���D�o@+ �BQ�Ĵ��E��9F7O%ʾ�+�!}�G���d12rΒ����YU9?T����I®</FWQ�)�"�q�rw �^h<ӆ��|�h��΄������gGH,����~��$YJ̒�r�]�ƯTۡ�0� c�yJ�K�(���fh1��U�e�F ܇~LG��%�$TS7_���~)��7Z����IJ��<�����iμ�WC�� ��� Y{`k���BW�1 ���V�WhY��:C	V�� [*�?�
�o$�a����R��xYוЙyy^�L���Ћ���N� `��G�z�òӇ*��J�ϣ��I:���}�;Qe��j�n���f�b��)I��<܎
��y݊	��B��!Ѧ+�:OGZ�ؕ���.,�c��Ş�4�[��|�k�� �)c�~=J�>�-�h�fG��XlxVHYEB    2f6f     ec0'�C�I)�m՜�$��:T�z�v�1n�����pd̲�<d�<Éldν��G~+��A�4��<�;4I���wF'yTL�w�4�0� �1��Dz8��{�Ӷ�:_�-'��lLH*K{(�:�vP�#\?#���\�G��<Y� �䐭@���P�O���ކ9��a 9 Hǘq<$@XG ���d�Gp�W��!w�@�f}k�[7#�.��5hm��Q����C���u*I��)i�ax}ԑ�P�#�@�'ea�G�֋�od�`��V�*EN+�����+�i0�q��}J=����5��+d�4=�z,�cL/"LQ��f�����K�D-*����i	�+W�w���&"!��ʘ�3�Iq��Dx���� �K0y�:sn�i�YG�A��<���+��rI���y}ړPR��yha�Gz_ڹ�ԯ��+���#~A��#@���s�cq�OB%c/a|ڝ�Ӹ~�z�#Ȍ������kB��
l���ؒ�����B�Jt�!� !�3
#4Y��4���Ҫ�	s(z�`O�,���.9�b��f����q|s�a�S[qb�F�,����4b�+ ��W.����r���nU��Y/��2l��� �=i!k�	����)�k�����;�-P�܌��<�)��Y%eg��N��6�荴}�gѵڪ���0�
��Ap����Ĝ�U�Ҋ�px�`��Q��7֨��m�&W���8%4�{��U&y�����U.Y�%��d�%�;`��+~P����i��@(u;����0Ŕ�KS�Қz��,�����@�:�l,S����^YD��ߟ�y��@.Y���v���Π�1J��x�#ny���s�`�F�����آ�7�]���>1�4�G��NI�sҾ�yO鯫����hR[4*�@���j�;��EK$����Ӛ#�*gʕ��XikH~\�u~0�5���"\,��"�U"��_�)�F��ő#*fk�,�4$���+��R��*<�sg�פ�O�a*���.��e��������z�:%&�P����V ����5K���@Ʀهe\{J�?r���0�\�آ�l�
������Mn��Ϯ�}g��nY���$?5]����ۦA�Y��Q.���Z��gx����Ε<� [���������ŔOG[jz����P�F=��+�;^��_�C�i訶N�����<��ȶ_��ZQ�Ս�H�_8m�P��]���d���)t�z�KHH=AW�R/�\U�w�@r}8G����>����(��gQ�:e''��h/?�x�)QZ��h1�μMs�ayv�!nQת$�=���֩�({t�G�z�����b�k��<¸�b�ee����_��G��F+����_'�pe�*֊q����Gq�t$Ȕ�TR��a��nqlZ�h��%��:�����Y�ĶH0®H �ӆ$1i��-h�܀�4��=w�&�%�o��P�bl���c6>|.���+5��U����Ѝx`k��%%���i��鿇i���ٷ�<���A����R����"�RF�⣔�@r��V>Y	�嬼�T.�]�LH^,�ď���1���ӛ+�/��R�G�|�f&I9v���;m�>:h���e�e>vk��R��}��`S��"�F1�;��d
���A�#h�
�&��|�|���>{}�n�h��y�`����R;��n�NVp���w�S�U�7�i����?�O�(4�`0'a�fϞ�dG2��1���n���ޮo����F>G2|�D�*�%��0BM�*&~9���}G�fz���a �M��^D�6�"��bkY��[ǧ�F������ �lzD���~��7n����)�1Km��윐��њ��W4�%s�*�"���x4���x�+�.#M�s�h�2V�vppFƺw����3�i٣CWZ,T�J��´�߄q0 �p�6��ß�b
�U��Z��\���8	5ڻ%�S�`
�������3V��n^��	���͇��=�� ��Z�a��%�lku��H\r�6��$����|��-3��ͺ�"I1R�zC3;{b�C���(
Kb�J0x�#Ĺ	�r��.ik�)�p��)(��vn���3���2���Xva3�Ħ� ��T@��ac�d *	T�	?��M�t ϑUY4�Iچ��3���r�#�������
:`�(s�8	�h[.��JmQc��p��7gj���A�����l<\��z�R@<�d��K~gX5�������	$h�S���)Z��2&����w�֝ǹ��Ǐ���VsB������H޵�T@ܞ��µA�7C-VsQ��+p��b5Shʒ4z��h��� �7R܂#�����]X ,��<:ߕ,xV�5;p nfy"�E��,����0�����B� �}T�a3	5ؒKT�[�s���b�m�<�L�⢻��)g�~���D��:.�s-�#c�t`71l_�5j`B�!`a�#��`͔tT��i�#X����6�D(~��,]���{��L�6�8Q�h�55W�WӨu9�뾮��ID�U����h��T�r:���o)��W�-��K[��bD!!ó�?2S��=d���m��@�!��n�����^CKz�p[iӔ��{�9<�-�����*����J���~S�����(�#��ljt�v�^-\��]č<�'���$�ǜ/n�g0���F�����`@7�C�&���uH\�3���k5��q��TTLS�m�P����:z0qݕ
�LWz:�Х,}��r��y���_��HD��������zQ��gC���)�	�߹���S`r�J(���X9�eH��$�V��g*1ʹq����rе�8��D2��q���ԧ��&�%b������ʗR �팻Lj��)���GU�%dV�g�}?�q1z��W_������1e/�X]��)�,&��&.v��K�P�) �q�A��V����fǃ��s��ʌ�K��+Tyx��ȳ�R���S�@2+�N�ݔ�)}ٮI��
Թ��u������)U�J�����*����i�=���5�l(�,ԌF���b�͖�����K�x�S�NlÄ~�YC�Cy����0��\��S ���٬mf#ⳮZ� 1���e@��(��[!�&�nj��av�N��~M�ː�N\�j��i��>`c�8NI[�NE8���{��q�*B8�J�8�T���$og���*{t�~�Ͼ�2�������r�W�YDظ'��7�"^[�)��ْ��0ݼ�wO��^���-3397v�PǏo����Q{<f�/E�"�ȣ#�U��:�ʗ�_Q�̹����8��J�XD#��9]��I�J��N�(:���G?9� r��R+n����>)��zXÍ��{�N����;��-4A�����ܰ��� ͹G��\�@l�~wtŇTARW��*_~�����EP՟��NZ=Л][���F�E�dt���ÀOٗ�Ea(�zܥy�א��˛�'H�9j�#�&�"d>jz��ˍ��/����f�dts?��L���n�.��m�dǍ���<���R�M�3`Ř弯����aӃ�%'����1L>���Zb����p���U!��Qcpj����N(��ߕ��"W�	I�VB_��9����M�/@���]�^"�`6���;�ǬM:��d7���������{�]��xBeOx