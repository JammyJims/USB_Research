XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����s������g2�G�A5��g8�/2�b�"������!aJM���kع�����I+ĝ�FM`l`2俇���x�Z�=ɎU{_��&[�������n�=�G�ň�mBv�{/w+��>CK�����pl���l�e��֠��lAqpFX�\�]��6#�?�΋g�kZ��ߓu�SAl��R���+m��&���'>�st�w���{��Я�6����Hk5��������<�(��NR/ܡ�W jL���n-#&Z�~��Q!�H/Q
����pV9�Zj�Gc��FK��Z�O�{�22��$�G����p�#��8�7[�UV��9�z�/�b����^;��5�t��Ses"libJ$%��W,q8 nY[��N���溣C�1>�.��8srs�Z#�BT�Bb��7$�O5�#���S�H�����ۂ:�����`7p�������옘
h�a[i($!�8HK���,oa�>������J9�X�vJ �c����;B�٩˞��Hb�ɇ���8;�c�Bɜ�^��$|���v��2���>����>h�q����������[�U��Qv��L�9)8v�88�e�B�k�$��_|�����u�Y�(�ap��x5���j.�j>������$X�QX6%���S%��hh�|10����l��A��
�U,�	�"c^>�>�;D�j�ǵ����c_'���`G�|��ξ�>f�Yh��+Bx`$��>�'(1���DyP�����!y�XlxVHYEB    1445     6e0��p0e�ҋ?���|1n?�_!��y�P�J�
�wfZ��#U�o�p-�������β�G��$�H�!�*;ɀ��gA,;���엾�~GQ��p�Q?t|�'�� B%ym�v��ӵ3���I6�;5�&���wYn�����m��`��{`������;��v��tLh2����s�UD4�نv>OB'�Q�_p=�e��,*��e~�~��QS�3J,9�(s�ܱ.9��0��$2�`Zhkx�޻i�+�Wە ;X�d��_ML_�1��BQ�T��)=�!�)m�K=���-�0��q8�e�R˽�kd�� {������g��
�Q�����@?�t�A�[�%/����h�	f0��ₙ��Ơ����-ox'�pg��Pӽ��z�V�.-�-#�*�l�x�BMH����h[�Թd߃Ee4�\nCp���"s���|�m#�˅y�Be��뗒�~���#�d)�B��x�����aqa�D?�9���ރW75%<֝����Og��(�cF��.��WW�E��G�37(X��.L��P�LpS��i�|Z��J�*]��V���6���Sb�
�[�v�.�����c�	��͖�LT���)�ۋ6�0������F�Ѣof��ϩ�$����(�a͞����,�]h�����%�K�a�D�W1���F��6ܺ��fI�V/~�s��<I=�d]E�����[@S_`�l��Q��Du��*���a�6�rq��>>WZ9:�c�(:��h%�F*r��&be�����bH�(��}� �G����E8�����?��NJ���.��-W@`���T�؇<�K���ƺ��DpD͜�;4G�~���K��c�}X*�{	[g#�� ���ŧ����uv�� ���6L..�*v6/k��\:�a%�~& Uu1��?�[qVqX���'��~��ų:�0*��np�����T��3��o����z[�gQ;9�QԖ�#��5�B��!���	ŠV �@�&#'���������V2��M��X��)��8w��k�Úu]�QN�vI{�.-H����Hr��~��|�Ӭ�+Z��T�����q쌘�3�OZ\>�	F�3<#bN�#��k��΄7��@\3�ҝ�jC�Y�w�~���p?wT��8`��咶X�� '�w��9�r$�$}0bͺ�WEcB��VQ�o�j���.���!��(/�p'!Z��'��e�v��Wa]9`�ܭ�#��$�����J������r�@+���ݲ�a�L.�s"��UaXF�����s�������0~�On��۽y3<<9N�������ھ�Ũ���Z T��`�M�n\��Y�h1e����E�޺-o�52�3a�_�J��8=�`�wg�ϴ�RG{�3q�=ٔ����zk�'޵P]t�+��?��Ҝk��7�D�?�!�\�BP���Y�D��ьF>XBJ蓺b����C�nPYc��	�^�|�5���_��\+��=B�f�NL��{6���;Ԡ�`��N`0D
�C�΃`�~�-��0�k�i�ұ�be�2�U��Kܷ)��Sr�
�؉�~qYͥ�DN��[X��R�����[(���M�S���:_7K��_���at�y���NM��Bk7��hd��:�D?���������3|�̤#�]�-�?J�?n�P�E]>^i&��9����Y�#�=.s�	�]IyP���;���Z��$�%���^�(���