XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����EȌ<���Q����k�nv�3Ȓ�VPKM?�q��LG�Eλ�U1�<)�p����\ܶb/94V���O�o2{WP�N�^ۏ���Y� �����,ǅ���t�`e����h9{B!G��Ī!�����t�æ�{`=���q�/Rm����lw�L4F()bn-����Ԁ8��s&�^ y�?��/)�T������y]o���g\`. ;����-r����w�.Ī�h��	�ïƏO���0� �tT{�W@b�����%/%U��*55jn�jI�b�G�m��]O+����
v8\���D��e��H��Y��*}���{�mݦu@��)��5���%X
���S��pݝ�C�x�}6�S����-�w�2�W��PV�]0��xbI#�H��e��Q��l��A�-52���7���WJ�3�!�����n TD�k����$�3���_p�q�5��Td�܆�Q\��0�.#�W��ѩB���G������j  !Ų(/���('&�!@8��s�e�o�FOF,�Vc���.�����{�[��$��f�k�]/�����o�[]�Q|+^{��.	?򥻐��n4F�uL3�8�=?U�vޮg7�t��~��Ul).�Q��3O���f�����_.|�	(�[aơ^��c��:��Ƞ�ͩ�]�vP~ī�Ռ|�{�h���V)��U妤U�*v6Z�R,�4Y�6�D
#x#�9qe�'����A��X�{|�]�U|ĵ��s4CKŭ�hXlxVHYEB    1e00     b20�%��j�Kyu�%�U�����Joo"
եދ���)D�ȕ
�B��ЮD���@[+<F�Ƒ��A[GP?��f_Y�q�����\ ����\�������`�C2s��ƣե�E��Q���G�Ӯ�I_8�������_lYhDF�~}p���E�`sDTP���߁Q�Ak	��U񚳶��	Q�
�)劦0�����@�������T�\l���5�(�$�.�qkڹ����@�{�mzZ���_�A��4�����DAЪ?�j_���0VE��M\�[��oS/y��x�)<�.��t�<�Zt`"T����}:�8J<�@�:b�;�{a��%k៱��4����!(t�/��h�F�.�o�X�r��t4�$�?�:1zd��g�7^�����`Հ������lIAY�c�PE��A��?�T���!���}f*���L�t�;��s��>�8Z��ed��@p�_���,S\�X�^w��PU v��=CؙP.�	��	MwV+�5!$�w#��{�o�B�`�R�}�"��Z;@m����W�Ѵ��y7�_�J�sȻ�=J�-��X�8ҫ��fF=./�qYk"��LS�+�$�����9�;�R�p���BR%��g�GDx���ѭ`@F�f�k	$!?�V{������y>t��'s�5�ğ�L�l�=,fߎ2�9��8�����羋'P����J��Þ!����qpE��~��N��[}\<�:5�P�t���IV(�S`���*�>-5� �ʯc��9B�~̇'^8� ��FWK���*����������s)�����DP���
�@�dG��[M���od�s�~�)?��"�E'�'
���
��r��a�`��Z p� R��q?�Ir��/��?��x�!���R�I�L��o�_0��6ׅ1a�'h'�6�N r��,Kw��CW%G�ҝ=��!�;l�JTܡ(C��R�i���r|��i������յVdo�
�6�zoL��X?��yc�_(�6 -�z*7� ���i		�G�`��/6T 6|CW˨�M��.x��_�p�H���'~���E��ʓ�66�J�C����,�ɁG<�t�R��w;d�j�Kl�X$����'���톫�D��n���l�HjY���AQ睛
�ڙE�2�&r�����f��gQ<�S����*�s�ϵ�ۻ��4�RW��.הa�g������M=D�AlފȞ3�������������&�է�f��
����̏q=��Ѵ�{���:�����jQ�#�ltn%�R���zYQ�*x{�qH��e��{��;&{j?d?*�t)wA��Z�nMx욢#0S&��=��d ��!u�w�8
O���e�n�bo-oqU��#)��p�[#���
�Y����^Y���&�j��E$��Z��o�#�q<6�;��QH�A��h�JԺ!q���!M�]l��6'�j��3��'qm��܋j���Q��+��]�RO��>��q�$�e��/�D�����+j/��xن�f3kH�)�V�MQ�ï���� �akZ���4�}����=)����J��F�^k5q��<4o�V�Y�/-D��� �����uo�(���J��	f@j��YB��&��k��.�:o����?���@��_q��c��
W�;�mʧ�s2��pe�H�Ǩќ���ݜ�f�[� ��e>�(4��SG_|<p���\�do%r��\�q��,
!,����c<h �Q���h�D��t���r?$?������[�%X*I�Tĕݣ^��s�!Z4��lpً�b/X�~��-�Y(=���l��w��1NXD���"z_�Π���y?	{�ڵ�+�?@3���!�tHE��87�45��������ֵ�`�!ȦT�D�����~tt��d1���-���ȏ⚐WR��l����$@��>�z�!�[�6�S}�;|������T[n�ˮ%�B��1��|��S2��L��*��	���o,�W��e���o�2�Kxmg i�����o�T�U��_��h9�0E_���2�Gw՚\���
���5s&��\��#�/>R�D�����v|����M{�L## մ�t���޸����K!H���g4��/L�Ӗ}��62m�^��cLg�.Ă��T�2��m8���\8�Ԛ�q��Rd�p�?O���ud���A�����s��E5�<��:���^��=Qh�z-5��hB~�$^8�/�o���4�*��6�!,��l)"�o��\�Aj����;��dϋ��\�>i��;���!s�����)^g�`e���oIΦ�I����M1o�x�.`����G���ܖ%��sC��]��!.�\b�=4������(�
N���LS���t�fLK���z�I֠���Sq��虜�جK"z��iJ!� �n鶬����
%&�9rгq(tdDڒ�F� �9��? )��ބ��o�n�P I���x1x��6�s8ڪ���WN��[ͣ�E���A���N3T� UH3Ю`���1��U���(��x�cGmt��-�����vm�;�y�n'�ꂐ��]S`c��5cs�!DU��L�az�,�
��=�F}�Ǐ�I��#�,��yQr��&��ɒjH�3����(f��<��D#��O(�j`(?�>P�5���������.nu�`ׇ7N�9�5�	�`o�%I'2��4��;�0��"�|�,�V�D\�� q���"���w-gO�����zI�K��Mx��a�\��%>���}�L6s�/c�N��d