XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��SE��� B� ��� ��-�d�
���+��t�\�V�I�dD�mMJ�ɒ$��->�w�+�Rd�U&(��z�K� �a��]#G�e�rT�ŊW� v�3���:�`���qm��n�'Qv@�X�2I<�s�����P�u�6�&��(�,j}�W�� �le�֓�Ȑ�/XӁ��O3��T��`�,~`�ϑ���Y��qEpVt�3}-����r���h�}g����c ��=�Y-k�Z��ϱ8t�~[��3�w��J2\j��g���Nx�2�����" �߹-��Էq!��,���4j�!�Ԑ��&�w-O�0������E���2���5�=���ЅC�M]CL���8D�^��&���AF�'�q�w\��N�$5�����h�V�8d��gg�LHFn{�i�j����^���~%�9Va�Kx�C��xi�_{m,`�˘S�]\����TB5���i��k9����rnO�������I�A����m��}����	�@�YQw�K[��K��������iO�3k�&/XB� ���Ft�)ռӛ������p�Q���u�a�%�뤓f�&)��-bJbp��� �84�5�VK}���oѡ�fkA�ܬ�w���%��[�g��_3����̈́�M:
�x���f�j������Z� �so����xD�lY<֜��P�gDc��~f���O_��Zq�e�=�6���;F/�X������^��y��)2IɈ�2�/PTO�l���N�uY�q8嘁� ����(l�XlxVHYEB    2aa9     e20 @]s#��T�OB:SwA����Ӊ-��Q�
THr�aD�����X>�ۆ�%��6�2��+n��� �y����͟c�K�؈�0�`�������9
W9[U���E��?{'�rJ�g!�K��e�B4��N�E�Z���#�-�"V:�g	�)S���#��\�ۆ�9 b�����}���)�b[�r��+�_z��o(�bJ K>	�C���&V?-�n���Ź��V-#E�\7�a���l�&��9 ������M1"d!/��w�$�]�Q� �@�I��`����s�/���Ȯx�3��M�m)�#͂�Z��lL�.L����Ѳ�m�fB�4".��+���~+>(:��<O̖���9��n�0%6~�n��˵j��5��=�ۙ8��~����U!�T d0t�і�C��g�(�) @0��+�U�&��$a�
^�����:�r[JOn%d"����Ѷ���I�N�F��޲W�l.3�D�n9�l��Ο�ǫ�U����ˌ����÷"�B��9\�^},�'�{E��J(�m��ϼG!��#�[��eQo3Y��f�UJD�J�W^�@��J�D^-3���ص���^�i���?^�w�w`�Q�b�'|a��Cʕ^�)�P,�
i�RC+�M�����r�[۫��FV����p�H4!3ա�6%{w%6��X��w���#8h3�)�8���5�kOX�~��g�O
M2����z$۪��ؐ��PϫT��g����K�8�,,���R~��:2�.���_"n�g�,��Vlr� ɣ1��K�]*�l�,�K�ʧ��a��_��ɱ�B9V�ԥ	*�g� ��n]�:�.D�;������6)o��4Oږ1:�/����A���M���U;X�t�Oy:�K�$���%�A��LI��� {��Y�Qņ����;}_G�eWf��4:!�z���:tMupi�:	x�/�)�9�_�c0	��`1q6Uo�~�:����h�a��B�Tl��G���`��T9Z�#?ȫ����Z7LOZd�B�2�oRרy<�W��E�4R6h	=S��"���n S�RW�{�T'Ǯ �1(Oԑ���s�8�ξ�|��5����>��J�U8����t8�,~�4�*OcF���kS�I�}�|ЙcT������0��+X�6 �/69$}owbFsa�-~�Ԟ�
��~��^%L6--N4Sl� t,��ސM�6D��,,� ��ű���4�h켠w�����*��$��\���0%�81B�g�:����^Z�� �j���X�d��|Gx�.�8H(�	b��!����t�u_�o9�1S6�(P
dp�#K�ieA�/R��Ym��8~¥��s���� ̃W*��4��x�w )P�9���nr"�����
��K���(�]�=���V�1��t��}"	�yi:���7.�D?*�y��[��M~̤�N�p�˄ﴛ���k%�q`�7����c���,p���5��?�Lߧ}�a�<�`���@�z��:I�FZ��#d�ꦹ	g�`\���
�8�C�9����Z}h�%��\���f{a�]E"�{g)����5�瘁�=�~���!�]Ǡ���p�����pa\JF��Bhj3s�ƴb��-$��Fް���FpO%�!'f�O�*Eg�s3|}\L�H���h`�i�̢G�dr8��V�4F�*�FY.�9X�Y���O^-s��<�	9����HTI�b~�[�|!���A.�y�Q?Q
U(�S8��Ϸx�wv�P��F;ӠL,����]Ƅd�|H50��O�7����:��x(\J y�� �P�*��	�I��Ҙ<V;g,�>��t��ɎrI��7��G��@c�!28C�p%y��m?��{�>OW1r�^�r��$������/)��/Rui�EP*�?�U0�<�S��HS._m�{؞#����?t�p�V�P%y�OM�,�O&���@�	"�	gU��E�8͟H�+��������������]��W��F���N@

�:g�J$q��@�>��/�
a|�wX��!����gldr>&��[%�7G����|~f�ǖ�`���F��;���XC-�T�?�dQM���JC�v����s���.��)�;�.6�RՆ1��4�5����'y��G:%�J̤�5L�m��!_C�����q'�����fw���ˡ�zih4��|��I{K��N����b���M`m������]E�kEeE&�D@��\�~m�y@�8n[���$wz+�r�wa�c0Ezd�5�(��b�1�sa��3/UH�Ȳ�揀���y|[K�h���g���{)�����W��\N�f��Ml�q��E�=F�4RI�",�N�2��þn�&w���S:Κ]�h����)��r���~�ԛ�99ݑ@��+�G�՘�AW��1����s��m��I�����F�����[UnP�Cnt2� �m�)�'�DQ�$T��;e3V�x*U�!���P���r�1�C&�5z�R;�e�X��/�s���_��#=6����-���ˉԞ?����1!6�!��1RO�d,,� ���=�f�V��5�Q���[�����-(NC�RfM�GB��!;�����Cy�-'�;�Q���W�5^�2Q�,ycte�@_$8YS>5���"��~$�@7\��H�=�gȲ:�NqfA"������68��v���h��׭��A��GH
�%�J�u:G���� ~�SH,��%P���}`V1h���`V,�7�3�g�^s`��R_��'�����w����K�z�bDٓ�И���Ti��"�!���'^�ɩ:&��>�:�S(��;~�P�m�]���ja/59D !f+��Mdp(a��ޔ�s�),����Ia[��Y�̀X�˵K�DG�P8'25ZA��D}��O8�9��Gz�}I��R�L�����,����^�"�<������������eG(�ժ�/�;���4zMs�y	��Ex�����	>����r�I����B�<I�.��\��96 �B��'����*�Y.Z�J��N��>�-��+�\�{4}��7��u|�袳�6�?�����`E��I~?D����^�)��������t�h�sI��-�5�=�P�������H�'�Wf($�۟��D~u�[�b����uU��
̠�x67q�79�feזV9�O~��}^X<Eo���-�B����Y�-�"���,��(�/��DMO����,~������fI�y,Ei�F�tvY6�`����2����9M�/����׬�KZ	�؃���>���s��S���"�2�<��cI�2����mgհP�����(˵�?W��V=����m�Z���r��w�iU'���T�-X}�#�\9V<�E�U�	�f�4�X�8�:׿K#�]-�P��̖P��>��x��1d��2���T��~����r5̸�6yz�E]��_�`�/28�s��;���G�|�?g"�v��uq~��v<h��� ����"��5���