XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C��%A��<kS���z	�+�՟0dCQ�U����!�yH���gv=r{ع�w��U�wS�C���rP��ބ%�W3����,xEsҰ�/N׈�	%L�e�ͅrj�
Q�]5#E�aΦ����V���&�y����H�}͂�*��<X?��։��,�t3.F�Fn3�6G����B��-�� �t��2쵳[Y�D�[����.��r�T�GIƈw�|���Q���qwK��:|q�# Y�*��ɜ��pF��_�,�f�"a�"���4��H� �зy[�й�Ǻ5s34K˖s`Ϸ@F���� P0}524ll�`V-����u1~��
�J3AR`�|��7D��馂���������8��4AEH��D�1J���?��jW9�݀s-@%m�Rsߣ��y_䪖̿�@��K�Cj�0h�����f:��W��s�K�5<�"����o��5�4��:L�޺m�t�����tet��)mz=ÊCf)�7��r��s��e`���ػ)��E�Z1��޳"�_���YJ��>>� �T#\<�
kO\
7f�&%�Z�`d���꼐�u�S�k��x�I�m�������e��٪|���)C1Deۙ�'�bOt�s���鹽fHr�|��m�*������2�e�6g�	-͈�-h�.n	$�����@��Kh�w��֤aό�܈T����"o�Sm��d�~�T��"�.᜘�P�U����h�1��E5ƀ�>��%�&���X@xy���B{Tcn���@=O�XlxVHYEB    61a5    14c0s��6�kLw��u��kwH�Xz�_C�B}�����D�N�T��n� �\<�CLu�hZK�7U�k��W{��t�c���SQ��c����J'�5"/pp�����9�&��S����N��B�e��<�>2sF������cP�*Z�3�W�1޻��+˓�@��|�ﳫ�9%w1�	s�˗�H;i+m_&��1��6�܉K-�j��6����`V�!�uT�u�A�tǋ/-�!�Yg!�����IyЏ�+x,�A ��g�$�1�`]+33�!`��8��͌Mы]kam��^�N��M)��b�qk8չO�|ub�?y�%/�c�����g�c�Z�&
+d��-7^!���p��`���C7Uj��4<�/G fl�|ζ_E:&x��w]0��}�ܑr���=8���`������h�Zw96�����uX��+�b�#L�z��x�Z�K'J���|`I����!,��ٸK�N1�C�U�,T�0jW��0*#ɑ�{S�]<��؛̚��b��+��+ ��p[�\.Z�� �y��0��+>�h���{����/K��(� ��(}=ܢ_� ��������꟡�TH/���vBm�����s�!:��%]����q�e8� '�j��D�j�l����3Y��	�:�#:��1<ļ��ͳ���`��i�I!��8��a���h�Ɍsm�Qr8� X�dm]"�q
2�4���-ސa"�x����'yd@���Tf�B�0Vx�Ƿ�p4��H�i�����9�T�"�$w���cTj3�i��xN��Q�/�W�\����J���y�S68�U1<e���{�_�'��m7�����_蹸J�+��)�Ƨ�1Gi[�j�E�R���b�o�a8�,�*�6 N[���ѽ	PWݓ���U�bY
^!�����5�m�����0�ȴ�H�o��\���a��/�vb^T(Sª��5&�i��~oeqBF��WdA�υ�����)��8=RS�ѨA$���X�K8�_�t���\'�����4C�z`T8�e�:K��_�^_	��P]������PK<*����M6j|���d򈬩B���䮜�+PU��'8䯔r�a�pwvD���:.�thS�)�fK�+�]�6�R+Zs~�@g��E�I��yҊLW��0L!!k ��"�<���8��9R��-�ŊS�2���A�=�?�)�N0�����k�=%^X������ ΊY)Tf9=}�@ ��.?P�
��ģMX")�VO8��J~����x��^��w�g��f��A��%�Å�o	����`l�7饰�d�-Dog���3�s
J8�p>�7�3���q�����⣖���S��?���Y�c��٠'��CB~���hΒ��=���X�Q�b��\�X�����A.���,�_0=�l�+bazq`Kv��r!�u�y�?�y�gd�_��'�r�Ch��f-_��*���_q.7�r:}R���R�7RB� ��f�g�>ʑ���|�����鸳��D��pXXlb�x1cKn�?Ë��k��1����$�Nƿ�\zh�K��.`Af��3ǹ欉M)H��B�( -�Q��`�v 1!5j=�s��
��'���=?���>m�5��}�,�o81$P���Ag oj�����ٖ�0j��g!V6�����$�\	R�QE774a�Hb]��ɟ���F��nJ�eKv�Q'+����й_YO����[�@�02��p}�c;�qa��J`�֢����̪F*8K�������,���] *��G[p��4������kF��1�UO���g �`�op�ĉ`��{���]���1�C䶧����U~U�����8�z�oP���86��{��RM�L3�^|��T�"�ն����4q�:��4n8`	�[���*�U�c+ϓ�>�C�w�,�i$��2��+�״PEng�_���{sw�B�s��j���5Y�U_	�c��%M�3��8���=��69��JȼQ���C$��Lo��h�a�Y���i��S���dx����?
u��ѡ�q`�CҜ}�/o����J�o�wy�]3����g�_��w�k�."(��3+����#M�^����b�Q����8�&����ɹr%���ç�����d0�C���Ps!Kݖ)ſ�Ek��j�]�w2U!bp�Ih�}�ſNqL��!Y�O��^�� }�c���i���K�T��b+v�z��2�^-����\��Q�z��~;l/�I\.��`��;J����}�z�G9���hﲾׅ�Pn ��I�t����|�(#�W�R[Q��X8^&l�}��-xz���?��]�p��*\,�n���7�͵�Nq�i	{�������Yt�Աǭ�q�Il14ʜ��&��?�q��O\J�C<�yQ�'����F0���^�W:����YZ��݉�l����!���!� �o#�
�^'��0h�=�:{�*-�ό��jL��= ��I��rb$2��(��M��p���;�"'Ӑ�U���m�A�&�g}V�]='W�B��8![�����ZD�(n�?�|H�!��}rYG���,�t��GV��˥B�*@#��l�;��_�K_��E=�j�;\�mY(55O�&�ز���n��nƇ�.S�')[������F�Z��➌n@\�c��:��tbhF�����W�I�+Uږ�����Wm��]��l�]��	�-�dy�ԟc		��l���M�qaW�I��y�?1
o
��0T!i�fa}Ǎ�En/IXW
r�N��ey���=��ub~���yI;9iv�#�����X�иo� c�sf�a�$�����ob+i�#��M$q�d�R�#_�k��H��u�D�CR�@�}�e��c/а�v`zze*�}���QI�N�g!�U0��l�h]=���̂+*�U�t��KS+BM�)w>�1T2�q���U:�w*=�!��	'�L�U%���4'w��I���gh����,V�be� ��<}��ij�麳	>/.��:��eA��$�/��	�����;���g��� ���d�O��>h_I�(���L�n��=�	<26�ܠ:�kb~�����+i�����n��%�	[ɜ�g�>Ɋ]��ݖ�p�f�e7�A�j�eX��`H�l���Dr�T���مNqx����1|��F�-x�\>��i?���Nu=�{e�ǽ=���<w��U�ng�����*�����I5i�Jd�bLBe�mM̭�)�=�.�X mm���kW�{�@&m����E4�4�8`׿�m0�E՗�V�7I�e�7�6���)��*��Q��W���D�����|�\PӿT��:�v�N�=��E���+5��$;퇯����=ky��3%��U^Jj[��&^��90ቝ,z�nm@�����jH*o�
{���?C���/���#UZWV�e/K����s�6�?J)�D�TG��ag� ��B�_�LPX<��e���B��Gj�3�E;���yp�}K�G��M"��˧f�A��i�έ�U���k�1�zmѤ;l᩟��Hj���w0�\m[&7�+�7�;�+:�E�C����7�5����������Ԃ�	se`��d���l��wy|U���8K��ss�҆P��ef�D,��uE����4�U�c��\�_m(�#�?��N��!OD�K����,����C���۹՘��]���u\y�_S����m�.b�(����RQa\����5~�ŠY$~�)�+�����%3�	׼�ނ�J�=�{���G�o"���q�x�}�{��YC�VU���-��Ǯ�����N ��Ax�=���b�nm���{��{�or��Z��9(�	i�L��W��I����sO �fS�%�˴l�X���}��"h/��O����mS<6�Y�֣٤���Jg,?���4ݣ�!!U���A!���l�}�^$����\�,,�s���p���[��������Ȃ��iI�f�j�������v�`D��i�e6��vR_ﹽ����wX�<ƛ���f�>��)i{U�zڵ�4�	�0`Ҋ=d�-JJy�~��8'!@=� ̗����O�wA��L����V�`.=�x]�X��QA�|b�,x&@�ʀD�A����k&i��X��
��6%�Oj�q� B�`�b���R(�6��a��"��?�-��B�Ai���$���$��!.� Z�ʵ���:֙O-�H9�~y���_})�2�P���ϵf�/���'��|�n�y5�\iڝ�����Rb[z�-�l��%�Tʡ�$�@�� �(5������oH�_t<����my�>���u+5�z�����0tx��z�ni1���k���MJئ_�[3�[���oȰ�Ϟ�x��
��v��߮�q1#��ߧ}� �؇��r�,AD�N����2: ���'������!��^0�Aw�_���UG�B�>/ԧ��}L	��f#��T+fb~�x�,�=�q����[TgI�0tSQMs��M �|�9�J��f���b!����ㄻ�W�]��eE���V[kA`9z+R�It�5tꮗS~�8D�KeᎦ�*j���/I^p��wc.�N��Mp=�ޟ8���m?}B��cG7	�^�^2F�a�K�!���5Z
�}����⷏p3����-�E��n�����v��%�Y����O7l �`����.�E��״5��$�����Ȍ��ƙg�3�/���6ۊjf��3�i���Փ��%�@&�R��+���wa.�=uQ�mr�}�)�,����c�|��qu5r�� ���X.���S�B��{L�u��G�	����!�1�5;l�/W��S�v���8P�C �� � mMxRn���]jDݼ@�#�:�(�W���Z��0�?4�M�����sŝ����.�x*�h�E�<tx�����'�b-qڐn��Z���1����J�a���B�!]� N��S�߮�X��üŧ*oAYHkz�'ǔ�����q���1���y�ɆQG/h6��V#�RI巭��(��d� �sz~����
�Wn�;�޹���0'.-�l#�l��y�`$BT��U��Ċ�Q�WS��ݠ{���s*�U�Z��\<��o�9�aM��'�ո�9������; o�X9�>�I��@�0�˨|�Pk�J�<�*�2���1��x���?wx��!����Q��A�