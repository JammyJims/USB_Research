XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4�t��!�a�KD�d�f�ʆ�,��ǩ-�-@;I8νN$��;�F�<+y�}ߒn�
<�;���1'hF4���=655tJ/qG�/?_n�q��'*({f��D��P1Jh���	A �Q�y���۩�B��L?�!YI �z�m���eCc��|sB#�v:��I@a[y���}�,�&�lo�0�-I��>Q�"ٷ�!��(�OX6X��iԜh_�k&�L���r�h|ϏE1f�9���?X��=}hj�J��(�#�gW�H�V%H��B��M��\�\~����T�e�e��X����r X(�O�KL���JZ'���ԋ�1���� ׈~v=�}��@�hg�?�I���B��Mǧ.�Q�����eI^w��Uϟ�k�iG[�mJ�`��1W������H��*��g����8������'ƪ������n%-?)�2ji�I��h��ģ�� ����AgY8QR���.�N$ԽV�o������$wU~ꎂ�R��H�)�{쉔6���k�ZJA�˻�]�_��J�R˾Q�/]���wo�q=�2vXzc�Jӵ��;H�:AǗRr�����?�5�~���D�=*�EebuЂj�r�C1[��\K��h�^��o��]���1�K�-�34U�����=e����� AQj|�����攉���m�W�*�:y5}�7���pf
��I�n}+��/ �]�BY$�V%�2�!��ڼK6N:�������h*n.XlxVHYEB    57f1    10c0.n�K3]���{q����,�|�6�?��Օ7�j�C� �J�is,zM�6��(�)@��Sc�������k����=��ܱ��F,aK�n�4�=7T#;f!�03$,�����O�J�`xH�
����FK/&���&�I�I�n�a=������ҙ��hO`�&jEQ��~ }�b��q%��B� ��#�u?����"z�P�?:�UwŤw ��S�Z��K6����T�fI�;u�<n�G��H�R����LV�����C�'����l�/�i�bD���sf�Wx�`k"v&Ֆ�k��4�~��y���	^G��~��F�Ǒ�p=Aq����#8���:��S���8#�|��\�~��ER�v&�T��R�y�i�e���=E	H��N|	���^���rswBZ�ͧ����X��r�Yrt4�p(�`k�6�%#cq�^��W�6�F�0�N���)g0&yPظQ�Ch&���W�^x$�����[v�'n㐍����gX��Fy-.ώ/~|��CK(:��6����>�M��ǻ��6c���r ��	R��mЀk��޾	Lzǲl�<���C�j�D���~���/S�rid��ջ�S�uM(�;����)�P�T:Ƣ���� �\姳������p�[^�t+wB�}t�Z}n�擡=3 7q<2«�;�� PҸ���sкѴ,T�fAwIr=d[��L_E��k�`^<��ڱ�����!.Շ`v��@i~)��Z��N�V�����o�?v����\O��jZ�:�T�-������Zd��F��ظUHO��S�N��>PC��/��\�ojO0���Y��A�'��O�F�B[�;�J��N��]�k�]�BXMJ�gK��1�5]Ï"I�a��z��UL��/o�NP�;�;J�z!�$���X���Q�Y)B�p�='�5X���-3�S!��l�i�6����w��i��|����1֞M i'P-t�N�3a�`$1�1a`�W�;vp���	�>��&J]�n���}����?��shp���"ߡ��q���ʬ@�ũ5N�T'>��D?����=,���c��+���� �#'�*
Yd&�V�Ar���]�k=轘�$¯$:�����r> λl���3��ـ��x�4�`e���"�Hz��864���Q�i_W�AU�'�@~)�g��K�ƚ�.I��O�%s�Qhd�KU�ZM�/�Д�i������:������4�a��7ǁ{�0�6��؇B�?.@�1>����>w��"D#b,�p�����4���AJo�_�t�AA*pmK�.5<����k�%�R�	�ZJ5������7��(��e�%Q�1���R%hx�_,���Ȓ-!i�F%^{�"2�+&)Z��g��
{��Cu{��:�S�x�m�b���S���7��5���Lp9"ۤ��_/��66�xoh��6�T�8���� ��p���7�2'�͇��	�E�-:h���ۖ�1Ct��u������NE%�CH6R�����.~����B��/���|)xѸb.�6oP2w����@��W'Tƨ���.3dF0~O���С~1��HE+dɼ}Cb�9�����K@���g&��*�����h��;v��ᵇ?�-aek���+�U����r��B���Ҕ�^g{��On]���.�@��J��T�8:��"���������KzH?<����2x��bq�=���N$]=9cxL:m��c��"=�tw��F���[��#�����8�M�t0� T�����c~wH}����Q0q��r�}A�Z�f�&R!�lF�%�u���3�1"t��D.4�|e�a��!�Mv��:�\��mQf�gIY]ιiIuoV���-g����ٽ�Q3��%Y�4s[D�#�ٓ�K�0�no��U��jil��/1��<V�������xe
B��T�����j�0@)GD�uH�
g��j�� �5$�'�2�C-��e��C���FA ����
 V`��0��П��,zЉ���H]�,\㻭	��҆�Xdb4��w܅�$�0&4/3.�:��V���D�����j��e�������D��Q�A�!:l�ɬ*�ƣߍ)�ܶs��@�:[+��<�Ҹ�s�B0���&�\�E���q��)������Ӳ`�'ҙ�?�i;b��U{�n��λ�a/2�j�r��P���h6�	�&�|ϋ�p\Q@�sF�#ګD� ��L��@�}Ifw�2'�1��D�`��-�9�*@��hL��F��+�^�o�Լ;�ˆ���_҅�T e)�+aV�� @�5�oV ��H���L�d��<��d��v?�����YZ	�^Q�T��{�_U8N�������q+Y\(�A�hy�g���5���\�8r7]��j��I����x�?)�Q�G؃5J�x�����$`t!]�!S3�o;��,�nuzˇw*o���f@�1C���}=���fi6���ߛ�����ƷC�c��X��{�/<np$6Z�����e����?z
o���0��m.Z۝5f�u���M�`��2yҜdR��o���c�
��wK�]� ǣb��7��	�����^�F�B�Ϳ�Xv֝U����Z|`ST�ڗ5r�w����`�Y�@�+(�<3�<Tލ�;O>!=��������d;�q�Xݍ�eӥ3�n����ĉ�DJ���z�=K�(�;��
�Q�=���I?Z�T�%��܌\� {v�܊��e�ڍȷ��wm��ܯ����eY �`!��ὓK���̘#��F��A�kO���@�"��\����<큫���D�pf�¢<�����k�_�ӵ��w�z�}0.�8H�����7�V��W�G);���S,b��(�+������FE[u��b*��l���ݡM�fP�/�c1)ϧ��j 󕴙%�sJ��W-��(-�f5Pkh�}k��������ţW�՜R��N�})�#t��Ԕ��ԁ/,}���4�$N�oe'�@V�ˋF}�
d���ec�;�±��<��| �=�E�BG|YO���$���ܴ�{b�ՇA��^�U�7��p�;�w��,
D{/��CF����. dV_|�.4�ރ@ӌ�������"�1<J��̾p��������i}��ε�H6@�f�_�[*�@w�o�aR���j�Y)G�Y���,�ܥx��7~Is���U!�9
�渫�6ؾ��+�s�������V|�ef�Xv�ٸ�x99��%F�I��pĉ��g�kꬨ(	?�k�tPRY�[��(]�a)�u���W|����h��x�Ά0x�����N䋶�.�����*����Q�<��j��r޵��5�*�U?��pa�e���J���}�O46�Ԥ���'�v_E;N<xU�V�����5!P;���xA]T^/f����K���^�r�\2��B�{kې��'1@��� ���o&h� ;+Fڨ�z��vr������ɀ��y ~�@x�[z�u���1�H/O��9��-+U�V�]�;��sj������B�G��<�T$9�O���6L"4���{A�E��^^Z��U�t�rz�P�X�5sT�&��F��޺��=Rc���TKp�n]�X�4��\	��4��7@�d�v��9�1��% ��8|��ٵΛy��w�%��	���gz��X�ƙ ��q��ݎ���m�Njxw��U���Wd�?� �D�]}F��M�&DR�yZv~�d�����W�o4'��(�LؿjEc̎��Ph��ɔer>�T@.���C�I�M���"%"��!{z��#���	yq .D�i18% ���v�x�l8Xa)Æ ��
H}[2�P\X�#�ع+8#"��&���`��>��}�J�S�X�EO�=����ȯ�ͮ��}�ňW�ht� �7B�������jr$y_�+X�Q��m�,b/q�{B��G����;�k���_��֙sѫ)�]����MC����^)��)�u�I�7R
�
N�S�r��M4�ZI�%�^a��.��s��G&̒m«���X�"Ε��U=Q[�+�6�`��Di�S�s|���-���9�`�ɸ��L�U��RZϕkhA'L)�4 "�����ɜ����qҋk�Ul�P�?��@C-q�Ti �
=u����4���Ql����!M��
��r�,�{A���:�gz�|�T�ڐ �tc�SЖ��