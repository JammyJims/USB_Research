XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��x]L��ùH5�NWf5��KnA;��эt8b~�	���	"�3���1E�$����N�9ڭ�զ��E|.;uk��y��,�:����kD��.'��iֹS%eZɾU��Y��0���(�f�O��5��L?x^�c�{���2j��a]Ȟ�D�����f`>s�DN7�E�&Y��L��Ș���*<�}T����25m\e�7�,�����JנDb��ҩ�U���¤�����ɬ{��kQەR�<��xL�P<n��e�1��w����m�|�O6��s�*-I6ŬC�z�r���L�ĢzD֗�	&�oV��\ҷcfw3z����V���kV��x`���9ɞ�Dᴪ���S`,�R��!��\&�=)��?���Z�0��Y����/U��N�"q4lb��l�jd=5���y|egk�Ɯ}6Q?�p�%xEb��(�����O� #D��ȟ���	@�渔���=�����Q�Jg�DK�E�����H�:�Ƒ5i�cE��SNT�6ﰴhݱ}4=���Fc�pp� ���4��Nu����\��tKX�·��y�e����HmS��k\��4�F�O9qM&����<�$#�^c���o��RvЌ3��Cȶ������<{c?=4򘀢��|��sD��7��!^��/;��2zq�9XY�FފP���E���,6��p��,��œφw�O^�� �]������k��!�6 xr��w<"Xy��4�	ǡ�� �wgXlxVHYEB    7994    1c80��q��X���xY�^YP ���\�^t�1�W*�T���֕q��aUUst
��� �.��K%7ԉ]����H5Hx���6B%�F1��|e[|95j��mBיr'\�������	q�Σ�&N��	t�z#�W'N�;uc+�LŘ�8K0�͚����Yә]m����S:[`{쩊R��-恌�.����H���M3�$0<��w��T��W14s�]�bһ~��5ʱ����g��P������BTҘ�Ԅ�"w�D��wP0���^�pm#k��̣����'��P=
�1<�#�-�]��[��jxf�#�S�V�ywA ��A�8�ߞP�_�q�D84��P$���$�a�?��C��hj�����/(Mi�D������#����"[��)�N�W�v�gU8:��:�D`'�i��	G$ ��K�+��r��$=�Yw�A5�D�p ����n���uӆΊ>��j��b�8��%���γS_NE��y��d*����sӬ6�է�JK�u�tQ��y3�$��W-��!�8�k����؃oMQ��!���:�}��Ĉ��R�WeJӃM��/������;I�V�p!~@��iΜ�Tر��S�� ���L�D��#����B��U����
���ѯ���_�*�l:�;b]��/8�x�R��=��13��g-�)L���Џ�}|%)��Y&7��|�5S���v�kb&8�����<wU�3p����0��/��1`%&�!�)M}����gbR��O��R�RZM�L�*�Z��LgN��H١y:p��gʏ2^�-���=�ۑ��h3%���
&���hM�ȣ1�<�gS�m#Je�͑q
�tS��h3��S���W��e�/Z������R]����bO�l����'�j[Ul�w�"�j�C��{3%/)[�:���c	O�!�������E�y�$Sh��B�g����#���Mc~A���5��SZ�f[��i��'�����N?��/�W ���,�"�#l���p(Z��W˷M�Y�GF8g[,�9�\SL��Tk;���!�'��젯�zUY[����C\�!����|����~")��O"�b��M"�Ï>1��MG��냷��am1�%��a㍂�NVQZr��1m}!h����e���$�������b�@�&<��噇(,^�=X� ɲS�B�����,��d����E�:G^?�>��V@/��*�/�^ /�Gt���3��I*��4��w�w��P!fh�����㛕+D�f�Ҿ�'�� w����摦9es���g|K��K�'}�����k��͚�T�ѯ��$jE�hb�i�%������Mb�*RC�P�*V�A9��]�#����#Z�CO�L��\��l^1Q�ʘ����bŻ5�h�'} �PY�V��1ܶly�m,.�&�4��KO��FhHlgV�~^���ap�h �����L�|Y��"��X�نYq/I�$;eTj����f���WN�	���5���0�0��(Ӆ'}zq��|�V��`:Q8�q�3xaNE�4���C�΋u��}��I �O���%q�'�{CXr�a�.Zfm�jd�̦������&;�nx�Nk4G'�M���N[���~L^�vܯ����@�9J@5�Fo�iI����f�c�4�UK��U��Ϧ�mWj~]��R�$�D� `@q���|1�Ԍ�vVk�Ŭ�y���t	?��RI� ��L*^fQ���Ƅ�XX������IG5���㕩����N��S�Z?@X��� ���a��	c��vkn0W��l��ʚ�5�����6�P1�5��b�rv�'Z�<�����k
�4Z�x?��;B݁R�p_�qf���W�=j�a�ND>����-<#�����w�G���s��>�,�W��H35%:�?���x�|j"�Z�<�np�ĸ&���
|�#j�n߄a�3�D/��~؎��˸)�`��5���Nc�y�r��r�Y�=Ly;���mo(��x�#�ы�޴!�$�oɭ'��_e1
Q�ꏾ���`��C�yp�'���ˆ�X ӡՙ�4g��9�Hu7��/����	Qkӗx%j)E�W0ϸ��5�z��x��*s�yͰ��sOf�'+n2ROz�X$�5�u�QB��{!��B��=��VC�-9����#@�BP�*	5� �%"ͭ/d��~�}u���ýA�e�0XKP�C��.���{���������h(����TB>
f��|/���8M߳ ��_�-L$a�H�����G��[5vl�`�������\��jL��^��$77xH1�u�}9.x�+��7�tI���"��@. �	o}'<*eJ�M�mD=��=��ӏ&��q�����mֈ��gN?;���&��?Yթ~jdz	��:���I��M'��t��
��-���&���N���6�5�q�40�`/z�X���pTr}��pw�|�`��fk�<v��S��kh�ޥ �1K�<��K'�o���Pw��啷؍�g�m��x6)��n�9�~�.&�������6e�r�!�n�o��>Y��v�W����:� ���N�(W��z�7��F���G[�2d�oŨWw�q�C��9x�a*�*\�\�k�⎲��>���?�Fo7�*y��c~&"P�7q�J�x�C�.��w��XG��X<�5dn��3�kP;tL~�� k�2L=���5;���(e�W��`�*p#kgC~1�FC���ax�va��F�;'o����_�U��7H�۾�|y.�t�[��\���`d8�����p4\n�P�P9��㗮u�[;�`�=&h�B���<�˃�q��ܧ��ɋ���P8�{��P�:7�~�-���#�V��'�ɩ����Hӌ/P�R_Tw��=u�k@P`}��\d�w��3�v�#xqe���v/gB��Q�2m5�LE�e�9�Ӈ�J�Gm28�����5ۓR�]��֍磌�o��Z������hі�gFp-�pϒ�~�.of��B��/�;�L>�W�"J*��wV��3�G�Or1��g�sq	��d��}��u0b�_S|�w�AQ��ٴ�7����S0��֊kJ������G�?��M!��*kܔr�q)�epN�LfJJ��Sk^�r<����Q�W�s�p��(܁87��� ?��Yi�	zF6��f���l���'룽��O�c�>���ajv'�$;�+�u�8���h�����5��NF�װ�f��1���Mo�Qh�(�4�s-��o������V�ͣ#�H�q����~5��V��w��z��@��� ��{5�n���ꂷ�R��#�OزD�!}�,KC'\r�-��z�^��g~�0�KQ���M�;�m<�n��U����sηQ'L�;�t�!�/����^�\JA����`�*e��ƹ�w.�X������8�	f���=](eB�󦺭&?���,$*��̬�fD��1Z'm�U%�*c6���C6���E��v��Nӈ��W�}6AtmYA���`��/a�eݔ�'����M`:,�S���' ��ٿe����k���Z�F,	�{S#���tG��V��������;��c�&!�K�=_F%��q�s��G^|��n:����cl7#��<�f$G� 	�n��K��BOh�����x�h�����Ô�aa��Xu:�zC�d��*�>�p��DP�	ԯ�d��v�&�oנ�1�6F�r�6\��O��Ϯ�H��*<HTE9p�N]Ms�����3�0/�>_�U�dQ��1�eX�(".h[�P���VCM�*ߑZDfez�\��"MT��B}���Aj$.
��=�0"d��+�+"�;����́D�\ƾ��l}:Z��E�K����پְ��&�-�fsg�!tW�,�׻WZ���B�	!� ��u���S��y,wf�gA�\�p��
��qץʌ`��f����2�$`ٳT��2�&�ޕ��������F|�Vr�<m�r<<�ˬ<)žѝ�7"����mҿ��&h�(�P�=lc��r�Tds�FL�g괯tv�g7eR������-e&�%�t����&�<�_wޯŮ��.ȓ��v0Cr�6n%Aiڰ�䒑g��8��gA_U"��S[*�r)�b`����^���n�/TC]c<`lco�T̋�a������c���=���3+S��Y��S!��]ĂQ��u�~*��0��N� �����ro$�H����4k�j�]�b�&]��7�R�^���Q��n	�Bugg$ӕr9�l^�D�]+��}g��=~<�t��E&4F�~�Nw�tsT<����~���5��lottn�`�n��c���w��X��.0#X��_�'�Y(��8)���`u���k�lBA��E)���=�gG�Hv�H�Y�����ܬ���Rr33�#�ڡ1��р�S�Py�E�<}��Io^)��Zw ��F��y/�]DJ�/���-Y�u��� �ɶ*����������������G����l{C�_�-�N�<.CO�ikJ��)�(�U���Q'#�g�CH_N��E�A�m�� Ɗ�TShT��wǃ~�ʌ�����ʎ�AbF�ϲ�mi��¦��ё�F�E���C@;>Ｙ�Pj�b�WU_�C��Tه���g�k%֟����v���c�{�W{m~j3���2����ܫQ�fPBJ]���1P��/��G.�>5�tԕ��2N�����xL�V&<+�;HE��|=1����'�͐�u@���!︧sn��s��BZ�k���V�ϩq�`�s�p3�-sR�O�&�jZHs�K���k��;��1R��Śf�Ei���)�n',9��0y�4��p����������ա@���Z����o�o��V�}v�!�����Ke
ܽ.��C���ء8s����%�F&M��V�.qN~�=�L��A<�.Ħ/����j� ��O@T�FTH�Nͅ����ߙ�L�H��"�A�Ea�60rKޫEJ���.���:�ж����Q��Y��m��.O�l�+��U%@b���oJ�D��e�襽������� ���!23����"��%A�Һ�x�/�"Nt�
����nr�b'��i4u4yCm��w�O�d�2��C�Y��l��݄1�t{L�+�5�<E����lgk�Hzi� �*a�2��LD��mIlt�Ħ*2��k����������\�C�����c���	����U��L��@+�����V)�:n)��'�d���o��
s�?������I��>~�jr��G�tμ$�����$N��0�3���t�Cq�d�>�p�U��N�4�bM�9Q������Ķ($��MF$�2f +�x�鈴�	LA�-M�9�o`E2�8��]<������V���k4 ���5�9�aS�Z��w�#��,ۖ*�hsǯ4���k��hQ���=�AN�@�s����vh�'�m~,t�_�`_T+�����n�&�T���l��� 8s Fx��& t��� *B�F
'Q�pwl,�|������{)j���u�ɀ�N�U�Y�7'��X�)\�� Cz�����BQ�O>CP;}¼(B�dԫ7�:<Y�7%��Oڙ���E��,#��t���o�dn�,iP3ۄ�rxk��6�
�I�7���*�G���hw��|#�� BУ&���m+�ۄ�����p�������\w��#I���<��� $����W{\#
.bQ�ێ���Np�}mN��Z�8�[��鋝ٙ��QA�Ai�Tk�8�0<��jG��5����uς�7�h�T�X�t��E��e�1�L�$1�	w���+l�����=c/��4v�����ĬK=��X�V�?�6
��VW_F�_TH;J��<q�V�m���)\�B��&�q�gm��`4.��R!8r	9�K�s����n˗զ?�V[�ԟ��b�UX��Zr^eS��_P_�7��){2,�;��p�@=:�!�y���xN�@��M�Ŀ1�#�{��'��/�v2#T�5�J�Jẃ�;GU�mB>N׈&fb�pn��*�:2A�]ne�����xI!�[o��� ���˔�CQ�!��`�1�S�� �Z޿���j����؎����߁]�p���Cd����o,�pq
B}�3�Y=���Q��C	�� ^a�C�i�q����  ������Ù� ����WwJ(tN�?9���O��b���TD����-�y��ȣ�`�/�Q���%���
<"���I��0'�8�6�e��m��RS{T���<��g�Q��ߛ0N��
��]���xz��U�ݖ ���"D-��+3Ψ='��_K���+�<�r�i�YN����O�WF�!���&`͙�%H�V�\�����@.�6�P�
�W�̇�"뽥	��|�q���<���O���t��[�:�l��9��s�r.1�^�w�5�E��h�7��R�2�P�V����r>b����9���D�?\!M���1�g"� �[�\W����GAG��ß���9�Gu�@g�j�^�~F�㞋*T�Zt���������?�C٬o�rK=�bc `��x����U܌#{��ـ�cN"ɒ
�>C�@��`MM/deD�mQ�b��-q���ma��U~�q�b��:)ҬϞ�څa�b��C�Y��ft��C���*���^��d�[���J��	s���.]�v�I�k3F�W��E��qZZޒ�B��ԲFV�L��PV@4��+dȍ�)��8��j*������3 b�֐` b�U��P""���N�z�ɚ`��6��k&]�A%,���������"z<8o�U(Z-�[rY���ŹNO�B��p�(���8m)O �~O�R��j�4�UGby�.>���H�����J�ƶ�붜l��Xe�>]�vJ�װ�@�䕶e;��!r�����TL�!8j&��+,�]�39���yD�qJi׊�|ʳ��=�&HQ���.��S��Ȋ�wN���,"f�x�8p������u�oj�Ke +�)O�`��4�N|X�y�U���Wg|���LʙUmX�u�~-����w�-K��M��-#bkZ�e���g�AhG�ǝ��~jQ��Ϧ1,?[aߓ��N7P������|���}�Ub�-����I2��ü~b��e�RXD�W��E�o��MU�L���eX��"��y]nO��s�ƶٕe��