XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{�|Z�g��X�ŉ����H�7mؓ��[]v�ͧW�L�9�7�%�ߔ<H��->c��M`w|0�Ү���F�a`��:�L:�B�G���Nc@�}��y��D�/�vƋ��e��O�n�Gy��F���31��I勢0��Tg&u�D�l]��61�1��*G
�w�����s���0�D��Ae����w�5i�9{��H�X�S�Uj��X�����b49E�@�"XL��V-i�!)m�3idv8[�a���Ύ�#�LQ��h��`�;d�!1���Ɗ)����1fpiV����vq#	���.�K��S~��'
;��%<�ݔ ���U	�Q4X����l�-ՠ{M�-�@�ܝŚ۫"�f�/?�.�Jo>���duE�P��~�"��*�:#�z�α�c���E�W�����3ί��rM�����J���HcJwS�#T*��BD`lcI�?������x�����7�z;�r�֫'"���o����]�Ȯ��p"'��m�8#�vx����z�J��ee�PSԭ�"�&��ߕ��������s�ؠ2�Zd0]W��������������\���3i�jԫ�ʘ(GD>ٿ�rB��KE�`ִ���d�D ����4�2��N^y��@u���5������h��r��is�t�Q���W��� h�M�V�$�1��7��<��CJ�Y��Ȱ�~�6hN��^4p�i�W�����U�h�y�'�o@x1F�ŧ�_���)y4�XlxVHYEB    b51e    1c70���2�ľu�oS��������:
NM�"x�ji�iϜ���Z���@0>�@�n$���*��X ��Ԅ��`�ۯ��v���A:|�ó�#}��^=��Xv�����c)���I���~6�9��1�J �h�-������;����Rۧ@��%4nr�0�H���aɕ@W,![�?��N���9�#������3;$�Y&���_�V��^�؎�_X��ٯ�9� O�+�XH�CuR��	\��j� ��_��!�S�NK]�xN ��}xwR����X�������6����䜚Xۡ�-ω���c��2ג�����'�dF��=h<���$�y�_[l�R��v�a��%.$�-d+�<0ГO��x���\J�Ns]=�O}s�wZ�vw*2g��1#�+?��]~r�IZ8��}C��H量�C��8�Xu�H	'�Xy��K�9E)P�ZWa5����#R�����l�]Y���6�����B帰�Ff��4��#�+��B?��9KSQ�����.��tw�A
љ��2^&	�~�SO�{���%��t�l�E�I�wjʭ~�i�]��	|�WT�9t�$���I����8I�/zJF8�����ڀ�D�p����l��Pe~)�Vz�xF�Mw�l��YE�������W&}�ͻ��,����u^oHI�.h�cٝ5 ��pF����T$�l"�03�|�:qi����D�Am͠��[�=;�ZD�+�񅏇��X�k��e��9z 80��-��P�1M��������V)��`)�γhݘ�G��o��
���F����PSf�c-n$���@����"�lx �m-{T^�Mk��=�9� 3�u�0m�4m*�ʸ��qkU��yl4�&<��*�e ��"XRd[�me��D�wPX��ח���\se�b���柑��-&��Q2;+��E��h�����ۿ��/2���"7�p��n�!��������G�Q�����y��R(�V�A����!����j0�zG��m�ؙ�M��1A��9/�9�5�FB�kwԀ�5�8`*2OI��]t��r��m�]-�T��.ݕ��{���r��	������� ����"�U�~�����	� ���^��ļ�RO1&��m*!{f��r݉�`�4An~�����vi��g��h�S�Y�ҕ�7- 8��?MhR3��r��v�܅p�ɞ�ߗb���k��X돛,|�8w��궕�UҔP�=�e2�H�,����Z���8{�3�ONq@n9x(H)�=P��C��їG��b��)3"��{��A����	�+�]{�*�WK�~e6�E�ᑔ��?�|�Rh%w\_�Y{���ʯ�Y���.O���((?�NWPe4�i(�Gn�n�x ��eS��l_-'��2�|G��	m���3,e�P[	O�dK|�����8�_=�i�gE̼��5՗�%[KlWŌ��T�둸�n a�Z-����0j@'�ΛM�	}Ɛ� �2�۶�\�n�r�gI�HiX��IA��0_�x�G���c�̨���&�vjR	{���E�0ߝR���|�3{Ġ5,�eJ/��	S� �����n=ɒ�� ����)�m���$:c�I�z�����y޳�����yc���`x� M��F	�%�m]QGmJ�:y�_��ȲW�SJU�Xlh�U�����n;r�+5e�TII�N�������J�y�okE�`�=�[�R_WE�Z8�T��?,�M�ŷ4��0
'T�Z7�~����B��2l+b�ߢ��y�����؝�����Խt|�}pF�Y
�k�={\px�]A�A(�,:s�enh%/Yqj�O𵒮A�$ݜGP~�����C��Ewע�%��uoҗ��̹T~�x�-~^Fm��fVލB������r��fK�W�,�u����2(]h��2�3�T *ݛ�̚T��/���n�һ�D� ��ό�Z{�^cBU�I]�`���񹶑0�L� Y_q �'�BT[����\FǄV8��r�Q���������C�nzN�o��\�*�>
C����A���Na����89+s~�ª�v~x�[�*;��ou�K�?�p�������? \h�C�O��X����M�	q~PN������$n��+D�Ϭ�o<֨�iP� @
��-g�3T9�N�U�V@O16��u㤜t�3��gBA�=�Z�����$1TW�i�Al�?�켑9Y"�:�]+�Pn�JI�<��v���C�͏6D��uM��Rs�c&��3YU/' �/�h�MVoC&�uHVQѓ�1�O{ґ�����-���E3:� ��r���v��1���{�d�}��-�8	�П;������3N0q���}5����p ���ua�h;� ������}F�9͚K26�(�Wﾋ��^[A�ϟ�gT}c����^����ϖ�|��J�f���x��+&�/�"$�g'�b�6��`"(������ѥ����I���dV^��%I�S�����R���ӗ�(r�<���ݴ��ޝH��{KW��ڷ��0����F����:���_s�ݜ���x+�	4�k`x���I��^�u����������T� ��9�	��j8^��-w���<� .m��v�6<�K������D�ˮ��Vіʲ����Pj��;�z���������&��oNRC
+iA�u�&	��z��F��C��]V^�)aX��ķ�E�z>Y�m�1������n�ӏ�"-���?�^��[�<��i)�/O���|����[A���,���:`(�9���q���~��dv�R�_��J���s�X�&:ဳ��o_�{�m��0EiE>�B�3��rl-�(R�K%�G��zF�M2Dd"�'f�A��W/��q�J\K��W\��m�m����4��^t���X|��� �6�n0j�Hz$�.��`j���|�m���ye�ɝ���x�f��;C�2j5��0��P���,Fho�n���7}��	,$���C#&lߤuI�ή��gխ���8���@�zmk+�}�s�ߙ��M�4fu�	��ڹ��{�ȬSue�K�
�=��]`��Ҙ|��X�D&���]惚 �æܲ�rԈHn�C��.���/�����byG����Ë��I��O�H�.s7�����HVE�%/[!��ʩM6:��LG���\ EV�#�������/ˊ��z�G,��ǡ�����1:���G�3�1��;��lO����m�����"J���A�V,5a�j��!���j�%��Ǎ��ѭ���d�)����QJ��ufVs�,�db��?�!�W@����^o3{m�5�OMW��re��[H�m�BmE/���a��ҴՕa�f�㣐�Hp��qW򘯮r�F-�	 � �vc!����ˍ�Ѷ�Υ�w�$�;�]����%�"���j�J
b�	���_����A5���X�)8�)�ήg�F�g,j~ߏ�e�ڗ�.u��DS���O���~�ڭ�R��v��2	���O�E��Y߲Qj�l����X�'��jS�d��՟��7]�z2��	�sCv���a�D�"�������?���0i��^ce>��H����*m
�ث#�<�UϽ=_�eҋ$JM��'���E�|l��.TcR�[�"���>|�|<�c�ZY��)|ٛ��X�@��c(4��qZ��y;;�g<��H���Q>4!�avZ�q��o�`]��L���(�p�7�9�:���&h,�7��qH� ��X5y�p��)�vז����g�Q�N�o4�^��\�	ѐJ��6���`��MKV�"Pp������x�����UG�&����
�g�Y�']�}vw��ӭaV�Q��|N������a��1ߧ����a�a�*gU�ӄ�bh��.��5�O�K�N��[���l������ƽ��P#�Ηސ���KN��@Ӝ����^F����ǲ��>,��#�즴	}/��T_ƿ$��wl3��d���K�@YW6IkB�8���1���-��a>R�h=	!�����?h�����-�W���-�J�Y1�Rk�<?6��C���F˒���5m�<�]O.89�S�y;�P��i�-s�XR���z՘'pj��+�%:����y�	c��,VӖ5���w<�7�+l��=�� �n�H��GԵ��6���7<���������t.H�X�BU�71���`��(Χ[���B2��@y��l)�2kyq����{�.f0-�^��C�����8=�V_�P�O@lW*7�B'#}V&�4t��ư*��7�8r�\Ͻ_���өi��&��~u;��p��4ª��j:m��zd��b���X`�d�VAi�;=a������22jM���Fė�S�?�Mt�g�N��h�Ϭ��ՐmR��G*�PS���)����4FS���]�����#^]�1KF(j��u�&���K�$#6�p�@2̏��2Tۯ"^��b���19���0���ٕϪ3���uw�N߾�$È�*�@#p� ��׊��f��ԆI�ۜ��_A�I�;G2=��u�%��Tw��K!ټ6f�^�pl��(Ϝ�츘����/ƀf�9�AwM[��*7?�8f����x�4����۠I��������kp���X����Ϟ������R"%fi�I���k���~��� �0�>#�J������[�ii,�gJ�B��^reWM��\��+c�V0&;6��v�i�%�a�H�G��س�i_��X�!��� �T�֖�d�J��A��+q"k�@WR�߿Aļl��#nqY���S5��rN�N������?��Z�IzTU0�tW�s�X�M����~��`:|E7}Oa�8O�o����L�{ Dw�ˆ`�]*%���M����)"���[��4��=т�WN7�DH*�mnƛ�3�^�U��B�.j�J�ZD���)��g�9X���P1w��5��m ���R/�`�8�/>X�^@[��!⎯��ɋ��l���XA	c���-7hT�t�������EԵї! 
Ͽo�5��2}h�C6�Jbq�D�4���q����+� [�$&(p��B&@�/��?�I�Ǿc�H�N�q��7Ku���]�F�q������!��Za�QA�Qe|�� g���薋A0��O�y�;��3"�Xמ�z}���r��<`1Y�/ Ӡ��Al��k_>�=�G�"�a��hVJ�HZ����kRU?X�I	"�'�x>�"�[�l�G-5�����!��Y�^��MN���*�H���t��q4��B'�w@�~eO'�LyZo�}�wÀ��x�}�{�v� [A!�q���x������uY�@i̲h���9eM�� �؁KFR���1��&~��W�uJ�݄S�]z"B��WX�t�P��X�k�V�j�X��w�?+i8�g%��m���Y�8�������uj$MrSzD���]޾'��p�	�4ph���/T-O�MG&�Cf_W%��ŧ}�}4�B��v�q�9�t�q*h����ꌪ�M)m�����8P9^��JC[$*D㢠������Nkkp[G��QV^��^�-P?����8��6蠭(�����6�z��K������v�ن��^�*-�T��u���#Y��H�ٛ�q#�j��aԅ0p\�z�Te뾈"z��a��C�M��4j0Z��Dhy��'��F�D��v��SȂZߜE <�?��BNG��R첝ݺ�˾�G�2S?�P!�����w�����eLU ��1f��� �Lu�l����i��ݍ*���!<��S|s�V<V�!�(5�m��MY�_2�R".[]A�_[�
�׫��.�(j:� x�p��x�Jl�"�K����!=�s�}~čq�B��<Oq����ܗ�[G��8�eL�"%��w�*)��|O��w,
c���h��MA��X�?�qq��vK�B�&y�T4�FNwRuĠ��0�]����iA��t��/u\0S58����M6��;��5�ZG3P+���u�h��w���ec��[�����(S�$�2�X}Xl�qLN
�jv��_X�j�I����(ç�!���A+�5M�щ�"O�6�?� k"���e�����^P�@���֖ �E�ͷ`�O���>�Q�)�]q�(�X\I��a<�^lN�͗�נ䬳m湪�*�B���tfӰ_w:m����#��ǖ�|�޸|�ܩW�`���G��,��� �<U�.8X+p(�����N(\�g�+]�}����y�5��"��W�����c^!4KD�bʧ1K�W'�T0��5s
���L������g����������|��&{�J,� 3����B*JvZуק�6�+�/d��6��+��X���c�_a;�gd\+���rԟ*c���n��Y5��E|�b�tԕ�J罏=���|1N���vm.3|��M�U��2��ҝb��VL�yag9��_���Gw?�~&��
���#����͖}�L���!�|��j,V��Q�Us0vS�s ��'ܚ�����h�S�9	������q��Z-l��Ы��:
k���'W�E��'�A�t��Nq{�5N�u�㸻l������:�.�#Y@��D� �7� ����2Xd�q�X�<�V�4W}P����H�_���Qe�����$H�ϲc��r|��e�������`9e�c��ٵȥH��Mߙ�J�f !؅G����5�R�oD@w��\4T�{?�:�� �.�\���-��&����Y��R���,\NP��[x��9�&AvT��nQ���?a
}�7��YB�X��1s�rU�$vF�����iя��/ ����BrЯl�4z\�ߏ%m�#M�^��F}�P�$��V.G�p,O��=�;�������V8�}�� �8�%��E}j�xQ�,FF� �4aC���D�F�λ����ӳ��|n$�Z�[Yrמ�G���'��X����7�G�	t���CN�p����d���LF<W-#L��^���� �lP?݂����M�lZ����(��s�L�(���1}o�!6 ��0Ȅs�c}�O���OH�M��?���v*����:�G��w�����ֵ����7�hڵ6���EJ��bN@��