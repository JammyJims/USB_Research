XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����T[^��.0L�*Je��s��⮁�6����p���4�Օ��E-�|���v@���9WU��| P���@��]-�4[��Ssf�#�?A����z��o�r��ک+I³�O)���$�a-v�:��q�4�+4�h�BYBC������&�;@b�)�]V������%S�P����
3�}N�{��~\�Ma	�<^�a!��)��Y�m�������Ia/4��b�+]��g��h!�pyg�v�(����S(vK+%8���'o������a��b�нE�X�h��hq�A�mTܴ�=V2���߫͡���4:�%��
����;�z����ek�i�KT�d;�9k��+4�3�4��F���a�@��'�Z�`}�\[0tBۇ2,�.y��S�X���;�o��xAh��>�v�;M<�8A̫�	(�=��4/@��ܠ� 
+��{��0���Ȓ�e˜0�>|�����{w��D�N���em�l6y|}@u������N�#`k�[�]�;C	3�6�Ð��~�(�񷱀<[ެ@��:&JMJ��.��:шl��緾�[X��U��^�s+��E��]XN�gLg|A��9si<v�!���[�{�cj�_����lԯ���:����z[�P)of=�O ��ć��
���bذ}�=4~@��MBg��-�ՓڏS�  L(���[m��ˬ�c�K��%�4�<�p�3�
�Ag���-�}�<<p( ,�zXlxVHYEB    e82b    2b20(#RK��u��<��jOܦ��F��|c� �����2�,+��C1G5<��i�
j:AK�S�`h |���R��'��d�s�/��BK}�R=jISf�>:[1��hgZT�Q
�uu{h�q$��(
���Y%�Y�Қ]{T}l��^��'�߷e|�LaR�ĴG\H�Mr*N��b�ó��S}77�[
 �H�B6��+�o�WB��E��R����L�����.��}���/r�>�ʢ��rEmVfL�w{A ��)�������������\?-�5s���W��'��~j� �oX[Ss��$U3���:�iu�T�u�!���0�V��.q���H��7V����%!���(�����=}Ɋ]X��~.�XX��z�T�*l����iJ��4����PS���s��� �-Ԕ~�g�R��1x3�n.7&s�vDZ*9IfϯyBm.�p�l&��Ǐ8�����-ֆ�Iʈ�����ؑiѲu�#�xhf ��O>�B�e�2�S�m2;�ۡ�,�����/,��T�������t��6��n�3��菱��NF2S�l�C� i���ط�播�5�*5�8|�� ��	X��^T�J����v�C�o�K(������̼X����1���x�����k�wJ��?����hܢ�E�u��6%�8�l;�=����U�r0.�n�;����{�JZ�x? :���D�T������Ĩ�H	�労�ƕÿw��%���&
��`ҜpL�"��>�z2�����^��q�'�<m0ǋP�1d�O6������v�U��WD�g>����c�5؅�|,?���?_�a�����Ny�o�+���l�	FkY)o D�7��R�)�T&���D]�j�:�"��A),���� �}�;��`�2��y������g�M��_v�Y����������k���T�(�x���2��K�ty'	r0��Q�:3f��@FQ�:�Q�YA	�:l������$��u �0岵�to:���+�=aD��rO�=�(Y6x]�+�]<w�ݑ=�`�L���� H�q,�i}�)���-��`yC�Ѫ�[��s�0{u!v�Q�H䯚e+ww�ID��$��v钑�ԓI���t. w{xf��礈]��s[4*ic�YTk�hM����
2T�w�����b���a�#$Hƶf�E&�\��Ʃ�Q�:ͼ�i�g�O������x�;؄�G�\�pt
���ݣ]:�	�ﲠGP�f�����}�{o.Q��k���׋6����R��Ղ9��Fwr@t�BFL��s�{|��k8zH�4~�i�O^�񭮙�i:k�t�8��*�`>��7�p�$9�h�i;lh�ωb޲9��׺kn���Z9X����cFC��䃨�nB�EF7���u�����hm%>�b�\^ q���p=l���ܳ	�E�O�aꜶ��<�b��dLi�0gc�����C���@�İ�#��mY$�j��8-�e�M�1�i��/�1���v
���ַasU`+�ʹ���z�p�#�w����	,٬�v����p����n���!d�Z��4�~~���E�b���(�x��8ޮ�Ӎ�O��q,A:�|��Z�2xۡ�o��)�R�Q���Bj�0�J���&�[�aCh������3�&x4:�z�v0L�(�٣��$��ct�k����C�?�`.�_�!	�ؔ}ۍHә8s�ʠ�58e^�h�rs=E�P-�b��]R]���ɵ�4�(*N�O�j}0g�6��B>��c��X}�\��Q# c�W��v��vd���~��e漻٧��Nb�}���\[�88e�V�������I��@ɧ�����M��)�.�+��T�,a�����r�^sհ �SL��b��)�I�Fb������Ȁz���G�Xk:|E���&���9QI����,7"��^�=b��s�I}R�I��G]B���آ�d�m�S?����b慸C�u�'͙�:�5~<jy�񆺊֓4���:�k���x�/"��<�X��r�x��r��t�_4�
3��nRF���s�9b��8��~��c��%��~�R�6飖|6�	����qa�1Pq����/Lk:��V��b�7��HR�pi�aX,�4�l�zW�'�WY$��+�B�/g�,�UZe4H�
��l�����Gb��@�a��(g����(�6/"|��챒Q�2x̃�x(p�%,=���O&� �.���yK��(b�ml+�������m�$�����CT�dy�rk�s9Uڧ�Օ�PlF�.6d�h��������N'*���DZ����r�nD��.����J��XL9����Z�]������f�T�S,�)����\����4����!t�m�?0iG���ҩ��~�*�~�Y!��l(6
:�hu�c��
n����)��D*�'ـ}���*"*=&`��YD�}�%��[���]�\�.�?��a�7�MO����A>�� k���':Ԣ mĵd�
3q��]�ʚ��9�<\m�y�
��������V�hhI�����w�+�(yۥ4�3r94��3��+5ٴ<���^**:�5�Ы�0�����E!��B��#����<��V��ܝ�ᮎsYׂk��ڀ�\y؞GVC�A6*J�b��[��%�q����+L��L��-@Ѡ���Qd���ˢ��� _��_�}0'!#9meP���xry��n(�E�L�{`W�EQ�٨���"�N"x���j¦%����c��EM� |"���$aB�3ł��u1`�km,��,[Sر"��B�~̼�P#^GidJ��Y3m>�ԘU%B�[d���f��,窜Y{���᩿�^lv����n�fQq�
����2xr�h�Kڛm��0n�]�޸�Yk�]�.S�ϖv�mñ�J=jlWc�/�����ޒaSg]bu�����;,@����-��fF�'�B�$��6{�_Ł�5Qd *���+�?�$���`/�r!(y���bX�:�_�f��?��A��/�Q��)�����[i��5?�a����G:-`c����\m�X�1�[z��̴;y,�z��W�d������_I,!���q<:3�����.m>v9�{T��:j]��̬ o�j�>�"�A�$�p�;�D��a�m��h��w�,�v� +-w��B�O�_��2=�Y�ꋣt��?H�ӏ�O�Q�?  v����n33�a	���>S�sdw��9�:�$�%C!,�'L�F�)�S�i�](�h	(�,nS�E�I��ۆR�a�"5��@ЅiH?�E��lՈD�{#���\��j���l,�Rn���4�~����J�>��爛�]���^��<הM`Ϭ�Md�������>N�U�����m3��!+3=k���wpB8_�Ah���ìj��~�A����nv�g�`#_��?L�` �:�������%��)�*�������54
�x��J����ܩ�w^���i�믺C��#3s��qw���O�C*�5gO/� u��3��T�\������Gz띞w�|EK@4}����=�#V�S"qq�@H7���mwl,[k�B1s�u�(Һ��3���U�ӃQ�m|��y�����i3�N ��ݟ�穃���"����R��@� ���X�� /��k��>⬣"ʥ�R��9:�f���J�5_g��x���g�3��Hz<���f�H����?�T-��B�b��W���v��}r��	�Kpo�`�d���ҋqz/��Q�h��IНt���AJg�j+������V�^��$�rk۹�����C�Z~"�l�ޙH���y�@�����zhF-)��������T����j���]�`\�@��&�,^:���4�Ȥf����H/	y�+��Tp�98�]=LD	e�����u����J��L��}
P�-
 �d^\~�T��I�50Y�_���O��N���'�[Q���U�'8�Z��Z?}r�u~�Q��H��m��K8)��Ā��
K��^B�5$ɴ4�Np���X��3D�+��S+�]��FdK�v�K�J��O��+s�b�w�m�|�}�Lˈ�f�N�Ō��<+ N���^L(�D����� 2�7�D`���;�e�S/�O"�������w~����N����z��"a�7A�ДV��]&�\QRr���m�@���+���ל}��I(J���wLɯ,<�J����9�:��LX?��l�ך���!]���y.4�)x��du	x���@��Y��o�|������D�s(w�89`����6K1��HE�sT���G|�4�Xb@@��~`���_;�So�������Q�EW��M�x'�T�k�!��f��ܾ���T��I���+erV�M�O����܄��V��0g7b���J�+N�_�֖܏g`.��6�<v�SӪ�*��,�%��Y0�A�k����G(oDsC�9V���VG��5�x�O��9���8'M��,�*�9���w��:���`��F�qN���R�0��ߒv�����f');lBʇy��(�*������˩|,d�t2Z��*+���@}�Q�e�_���~xm��8�ǳO%)��E᤿=�(w�T�䓱�?��u(j��ptd�#���s����x���_C8�P��F��c>`��qDI~c1�[��|�v����#j�8UE���E;|�;N&�3q�nG9n-}�G��F/h� ����@��]}JDC2`Ǒ�=\-w^h�<�P�lr�w�#�#M9le�5_���ו�q���+/��C������t}o��K@i��Wcv"��/a^M�fմ�� ���t���b%,KN�`W$�ـfdW�Q�ZJs��S���ו+ۯ�|,�����2#_vL�+���"zJ��a�R��G���6 �HgOr�;�5���ǋ�z|�?�<qH����r��oOi�p�<���1��Ikw8sK~;ʌ'��d�%�ن[5j�tt`/<O(25tcI�oF5H4��V/��L��xC��@�>�>�_IH27�;!����K ��3Y�8]C�ΨdN�u�kg��V�2<�#y�n�Nf�$����s��2��C"��(���&n"S�n��Z�3x�c�	��A��s �0�4�7�i�� @�?T�/��y��|�����;F��<��9�Y�͒Ԫ]0m<a�"�&���N	����h��Ƚ��e�
;�NT�+�Cq�:�h�%>m�o���@Bv�:-���]��f>[AT]�	�GG��gΙp'�aY� ��=B�2ϋ�	$���l�n�$�ǳ��|2�{��/��`��;��^j;�K.λ	�����Ie1��G1K��tgI��[oì�f[N4��J���� �2%7}���G	s�n�/gow��O�������j�7�ZA��&������U�x����unx���׿�7C
�ẜ����A��.�I���S��;w��|R�0��������aN��o�i���B����CW��⫗tÚ� �;����VW���T1�yM�6��?:h-��7�r��m�N3��.���YT+�e�'
Z��ql��o�(��IcР���n�m����4m��I{��J��1�z��lXt���I��[#��^�zt��Д�}$`�y�������Z���a�Q$^���F	g���9̗����k�e���m�Ȟ���4��j�������B;�Ac�n�k��1�J�\l��慿J�v-�u�ɍ�r툤��=I��q#�eE�-�BR:>bq�[8�B��av��&-�����U� �bݦ��(�_a~nE0�<N�+�q��\� �����r�iYކ����!Y��� �n�S��:Q�Q�s�L"��N4���� ��>���iN#���7s�r2œe�yO�.� (4lP��AL��H����5I����TN���	�~8���T0�'x�vgە)���1�\������#�O�i<����A)&|er��l`�����b�Pb�,�������|V�{K����g�04���IP|���-ݿ:]�q��=�^
���p�%��9�y:j�EHk�F�cY�����O_�mۍ�n^:A���:���?��f���#��ٹs��}�Ӌ�6"n�|����NSPl,��l�Obh��A� �I��4
�����5x�������G����x�����
��؁�/tyx��FkB�]8��0dø����O�$:!��?:4�~+�>�)�m/�A���U�����d���!1��VS�=]��O���)��j-���K��R��_�]�?�Z��c%UC�`�����=@ԇֺ��.�$Y=
\��������+�3��{d�(�ߢ\K�nY\ ۻ�9�oξo3(��O1������4�o>Y�Ob�3��d�&��k�b�d���h_IK�j���:7�JA �]O�BY�\�2��>��[�����Z�I������l]��K�P�#H2N��xstU+ز���x}��'y��l�J0h�M�L�w��n�A�żxC��c�C�Q���Z�k��c���]�Pxnp���K��
o��Gj��F"�K��M�+{��4��	��3����A6"!���J;r��W�v�O]�6��{֮�a��r#������}��p��v ?	O�u����%���U�-H#Q��K8�t(��ık3�;zy�W�-����O���'b!	Hxu҄�hY>�7W4�y͙U��-+r��n��w��8+n�v&;�B�]�J��U��+��6�oF��%e��R�xa�"x�N��}���J%C`1��"���H"?�5�z�
�W��Hz7@��3sSc�+0/�y�?я�H����gWl+h�D�A�4�ΜJ�uS�x��_n��`<C�����ߊ��Ŭ=����7�晒������8�Φ$�!�.#<T��B&�y�X=��, �̥}�G�c�~�`�	A;�?��~ �7�)���M��Q7�&ڊ�=�%*^ͧ�aTOWq�v_Ǆ�+?	~2؜�id�4 6ks�t���^��Y�!S�h�������$�#~q%����˴c^��S�V?諌t���}�^`Xt(	}g1NǤ��g��w�:�Gv��k�޲øA>����2a�o�� ����X-5>��,L�l_�2���Y��f�TKv�F�Ѐ��Ӗ���y�z��"m�ڔr2M �4��%G�!���r���]��F��z���l�[�_����q>!���Ce��/bC��tFm_���˳����J<���"d��Q/gW?8�22�,Z5���YN9�D(����go�u�T���E��uy�ZC�
^Os7^�a�e��eY��y:1(����o|�T_�J���v���$�u�c�z�^eTj4�s�26x/l=�PH��Ӧ(t8̞�`����M��LV݃0u�׵*������!h��o���O��T�]�����i���$����[�.�e�n���
���3SE�a(>�@�ɏLٚ5 ���m^�Z���\���1��>?�nM�$�#��]�c��.�B�/��Z�d�y��"��v�p&�p��c����g�7d%K�5;I���"gj^�fM��D�(� �C���Ɖ����L�"����dEH{Z��4r�Լ� ��a����I]�-�2�U�Q�7�����5qsaz�5�H�6v�a��	���C7'�阣$a���K�J9o�(R�nG�%����g"��֕yY7��Zu;��ϼ$s�?��d�J�`��]��C�Ƽw�M=��\�U�%*��}�O�R�M�4+�L�:�䒨'}���;�8G��!��9�ũ\�P��ƁK�6�u±j֞m/L�H���oW$A�������2����k,�t�ٲ����Ǫ�J�5�;F�(�e�"�X���od������t\L�(VĉY�N��J�T�O��H�)�ɩ���o��WĻX$���5p�2`p=�$���?��Z� n3d��}�y+W��*M$�hvm鵦Y�}�dA:�ad�3'�9�AցJ�r���k����"0Ri�=�:w�` G�H�0Vb��x~_~��t��	�gj@Dޢu�V5.§4ǰ��Y@t�O|R@�D�����b=�˃�ܖ�-r(���_��ɨ_DX��~iA��JR?˝K�PZ����t�T���.&%k����6i�"��JÐ[Xm%�?θ�2�K>3z���8~{jN��*�{Y^TV��wљĢ��ltV��f뜭�D	SJh����Yb蹴_�w>͊��5��1lWFZ)�"�Q�1F 7�h�`���!>��e놺{;�²�0C�EJ�4їel�&��*Č.�ž�A��w�P'}Ne��޸�Ix @{��+C�#��䇃wBy�j%K9u �4(v��鎵��l4�{�#˝�c}N{�,ܵC���v��H���b ��;��D2G��MA������ޞ�j����5]ܨ�,q�笖�h�Q�e��B s;���W�8I�@��[�O�����u�E�|�]f�Δ.W>͹+����z6���O�8�կH��K�B�S��V�o��~�S�[3���)m�X��������Q��3���L�(]�e��VH�g9��--J�.;�����i�*�`=�t�:��,��`Go\��;�
�-����9����j~*�n��MO�pm�Z	��xf�&g�Ϋ��� l��^&��AM��7칣�������]kꒇ���<���Ǽ���X�*Y��%����e�p�c<��
�5�:��Ꜥ�&�����uKߘ=`�
�������]���E�\���;� �a�Z��0�R� �6�b0�	�<2|�G�h��ݙ�i@;luF�u#^�uT��z�*�q�������϶�]�l��2��)ے�wAϿ���f A�B�?�l.FTGaNԝ҅�oa�� ���������.�ф�n�,�g�B�an>�:��2ϓK��T���A�4�M$�[��X��kQn"�8m��h{3��{fI>I�Z��c��?�!L)&��������f����`?Dk�ZC"4P�i���@�׃�tM?1c��X�DFJ�|ܐ�F��#��H�o�%�M�d���o��{BM��qɺ#���o��Z]�JQoS����ϭ����/wd�H�U$ǚ�_��乊���DM�r��9�ۡNO8W��>�f�	R�X�����SB)�x-m`�%�y���SE� !�wV�bB�0�KZ,Z�'Y�蓓��+��9p͇��L̡ly�c�)�s�a��"��W"ˡY ��.>ɤ��c�4;�^��_��B�/��}�Y��K�5������p��t�d�C}���vB�J��x	Ԍ�z�#N�>ռ�"Sk�Xe|���FF����P
�5C�}�WOA��!����f�o��Q��c�Ԉ1P��/�Q���Qs�AE�%A��2���ucE��D���-�Y>HX0���f���qg�ߧ��\��ȸ��a�`��	!�����9�5��&Ǘ����1���OQ�dT��d�<L{ T3��٧h�r
�)�2,���s���G��{�IC�J¿��}���y�bd�Z���Jq�0�Art�
���%�����՚x%�]d�_� ��o�e9z9��5�[b��(���Y�@�p�yݮ��Dd|p2Jˣ�Qq��w�q��*��_9��;�R�u�d~�j�e?��E�s�a�Rl�p �0VX�uD��s���$ŵ��a��ԙ`��4�����&��0ZS��
�,K�� ����v�p�A04%A�eF��T{N��L��s����Q�<�.�m�na�G�'��v�� =���H�b�K��"�8L�V��������͍V�z?�lW���\S�wل�E��*T����ơ��y�h_���_Q�Zk-5�0	�r�LB��C��P⟔H��&��kn�oؚPE�U�!Ԃ=V�!��uX��шy��b�7�+��:r�v:���B_}����SG�k�L�!nU���!/ZF�l!̪����*/ӊ$5�So�Tt?���J�h��u� �u�xu���<�9+cEf��v��ʡ�2f,@�<�������,�9> �^�&�g�:�P������L�lf�F�j�G姼aX��Gz���awk��a��ԧp��O8�L�q!���]�	���o.�ϖ��y���R��¯�n�
b���Ƈ����e���i��:�4"��< ��ds�x�Jw�%��Kv9�1�r�I�yK��<:�ޫl+�5��z_�����G՜�h�xz_A��o�e?�.ُ@0~f�;vt$�cd�$�M|r�ӈ�i��R�6���X����[�sD_�(��P�AN��E� ꐱ�ja*�}��#����N�%(�����z�>��p�\�p�po��f��^��Y��ԜP�
�嘠o�\�y�~�38�. �dv�l�);`����/���)b�B ?�0�����/��ygЊ�T��~����+�hV]ܑ�Hn��f�]#�H��L�m-0 -�P�Z�y��ظX�_��Q��i�#�y�B:��/4g�? �^�Gk��ˇgl�q�g���xm�م�\���f��)_��T��CL*�Z��x�Q��vG�f<�8�	�P\��n�"��ҙ~[T3���-~������ β�NfU
��5�"tۂ.�8R�ԶטM��$�G�mک]/�ʚ��S���B��k�����Y`�0�)��3dHdOЮA	D��L��Q<��������2�