XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����u�X���}��1/Nroa��Mm>m4��K�h����Y�P}���r/�sZ�N����yq
�V�,�3~b#o���xD��G��ɫMZ�G�"B��4����	�S�ꘝ{si*�2(�Wgʐ��!.�u�U�z����R�� ��|��o��9���'}�.丹�P�1�zg�u�tI�����g�X� /S��\iˉ�B2����d��վ&�S�y�h�����юG�J��p�:������	���;į��!��~b��������M7��h��U�R�����։���ޏ f����C���ză;�3?��W�E��L��f�>�ۚC4,=�D@�n�P|��:!�Ec��:�&C���+Y
	b�����W?׺�>��z���EQq�w���2(U@�0/).Wz\��.ub^��"�	��|�I�r~�S�ɽAqk��e��S+E��V�����	����@�3Y���Z&R�s6�-�%��k��RJU�¿��9���x������Y�5P}��_jm����Rf��*=] ������V�:�����j-����	M����:��@��Nk6��!�VU��W�cv���
����
V|,�P���S�'����o}GO�<4p�/���
�k��D���~�ы���>U�d���f8H5��IX���s��/�Z�"�&.�쉶���Nx�,':�lǰ���b72�l�W������7ӛG�u�~�RS��˧�T��XlxVHYEB    5dde    1700e�:������~���9���V��-����p�_��-	,^B�x0��c�=���P� #(��Ɠ�#��i/2�n��B��6p,t��\��c����U���+x�$~���8z!��G*�U�1�ͮS���)�닊@��6�T�`�T�j}��6V��&x����}]����iPW3��s��_"՛�ņZ�ge��f�)�J~PK�q ��N�X��l3�v出߅�d��L@� �B�(�ٓF��.SN��>�gw2+�� >D|C7s9��X#a�f&k��t�v%@h�@8)i���f;e7��T�YԎ�Tg���Ӫ�SqM>.;z�iM�������}���V}���w�AW�Ƈ^cVg�J�o������3��U�5�4��f�Ҡ�7�;�`Eɠ��R��}�"�O�����%�6%�F�t�d%����P��n-��hzC�ݰ$Ί�w�ה�=r:M��讆6�l�|oWT��-$�A�J|�>�Y<�C.^9S���mcwx;*NM��A'���|��W Bd�f�E��aY0� Y/+ݵ�n�+rN�u�w.�57��i�C�h����y�s"�볲^�)��U��={T�J��+1��xf�1�+^"G��aZJ���P�ፇ;�*VF�yυ?�PU$<��ڏ2���������]R�>�_�{d)�B9�'���0}j�_D�y���dJl�ݦ��_�jP���-�1^7
��%Օ�m��W�5�f[�9%����R7Ӿ|c Й��*2eG�Ͻ�B@o Yy�5~�����:�`��l؉��w70@�=��o&j���s�a	�����h׭��� kj����Iai��\"�p6+�9�`��s
*���.�Q3XHv�n�ݤ�� ����e����	T��bVʚ��(C�(�cƨ$*U窵b�wCU�Z���G�3���x�/�h�.�x��y���?FH�	��$�|F�ڥdE#�a���-��nIa(D'�'���f�8����i1l���HeE "?��_.Ȍ�Q1�]+�Z'G����5G�@�w�x!$���:L��6�{/]��* �^qp�a�� 5�஁c$1#���P=��v��V03C�I6����RP?�� �����@�BQ=y%��
���A�I�xK�t��`[;�u��� >�0�yb]u�����Z��3\ݨdi���ݼ�#痩oܟ� ���Jf1���{��i&����(ɇ���}����������|��b��~�u����W��+u�o�<kꎈ��g��V�R)I3;q�x��<����M
}P�����b�h��=kp��!Q�]�2>�������ʗ���Е�E�l��o�k�\�
�}鼻/��^ۺ�~�E3ԙ���O!��M�7�JW�=���<���B@>Y������鶱����y���zWڳ�a�d �"@��8�1W���x������L�6۲U-����`�_?��-P?*�Nr�^�^��h9OwZ�
�-�h����x���VY0�&>�Qۃ���j��Xpų��AH`�u��u������voN�!�64ʤγ���y��Jʆ��&fѳ�^��ӫDGh����h@4�y"[笭���B��R���)#�qC"?؟=9n�,S��?B�Iަ�/a����)��`��	S�q�lg�����Wd�����/^?���d��;�і��/A���SHo�Ju�W���Óz� /3�I��g�!&jr)���Gzf�JD���sx�ʪ�h#�+�2�x�Pwd'+���XhHۀo���vx��) x��^ �K��*�P�5�e�z����=�-������(0}wa	�s�k�ȇzr�_�����E����aO"8���Cu��D͈��%�Xe
>�f� ��y^s���"m=&nq��S�=�¶����^�*���qq}�'��[G��dZ������3`����.���ޗ������)�����J��k��%O�̼������E�ż�a�~,Ea�8�k�h�xt};�{XȻ]���C��x��s[�o��b�l�����E��V25�0QA[��{n����D��߁�Y�W�lH���-�ݘ�/Gm���BC�T):C,$c��e`�w�
�[)�n�0��C3mi1�� 2Ƣ�B^:����Vƽcq�.��h\�[_v�Vm�Dh�L��B�Tہ�D�5�m%O$Ψ�N/�����

.�	'������Y,\��>YA}t�ĕ�#���PW\\�K���}��kO@���#����X��B#��2L�[��Fc|"Ɉ�8����(J��I����U�l>��2���dX$"Y�Qn���)&���[E=���-,4H  =��������tm�8en@���L��j�l7gI��lix�W�%�K�a�.����M��Pn݈)W�?��A����F��_��3�y�X����-@ҳ(zڝ�H���ސ���f#'R1=����� @/p�v�����e/P�tx+O<�`.ʍ@y3�Z���1����Zς��j��g���*���+v���i�I�qf�=��g^�릨�r�0.��0�гZ�]����GpO����GQ�&��Ӈ?�,�Y�N��n�z���b�|���{�q;��;��/� '��D��_40ƚN��(�����^U�F�/P�Rz����:��d���CbT��X+��n�x���Aߔ����A��?PU�����+�7�8���P3�2G�m;��Mn�r��qX(�bi��g�]�$�߿�^���1�����B�C���v�Ӥ�-�0Ӫ^%��f�d;��Լ�ia�Ic�9F9J=z�H$F�_c�t�{����\#p":��D�&�XS�B���G,���"��gf��W��w�g��"CP���]ɢ	eP`y���a:
�}�q�F
�	�\�r�M��xט/��q��Mt�I��-ͦ
g���!��yԫ%#����Y��%34nv���u��GEr@$]_8�R�La�5�M�eS�pҘ��t���}e����[
Xm���KV�"���4ez�I�_���سA��J3�j��/���P`��s=KB��"��
Y�O�Ҍ1��X�R�R��r��1�?�;�����2��FN��[�B�:�7����CX.oKq~$ҽ��Ko����r��	v�)�$�/j6�1���+�3�+:
U:�ĩ��,c��M"<�@�K[�V?��5���Y���������^�V�p���u��"�ve|y����iM�`8�.�_�#�i�S0��.�8�r[�j"�FU��\�73��-]�yvw�ᱜ���Wk�R����,g�`��<¯���)�%�+�����f{�1�v�O��lI���-E0Qt'stl�+�tQ�.��Bݽ�z��
D��|g W��$t��v�ZhT���m-�w�Ǝe��f�?N77fT�=�F:&��l����=	Yy�K^^�%<g"?4�@����F&bpu5�IᎲ8N���䎈�����,֪h���/�ݺ	�W�i�h��"��%�D������3�̊C�ᗮXZ\���'*l�>��8�����3�Le&u+�M��K��E��bAޏ��&��(����~�1Z.a+������7��E��Qr�iI!��|���Fg���t4s��Fs`�\��-s���S�C�
�YF�S��T�C��\i|��w����I����],�(���ܚ��z�g �j�v���l�	6 ��R�ԏ4�\B�o\Ʊz�x̦��hT?�Y-ZA8�p�q)��*&&ݟ�Ah��W���S3vƹ�yҮ����I�;+K4R��uv��ZU���m���s�q| ����y���VB_��g��ak�˚as�Z�ҁ��Կ�36a땘�n��l:��-FM"�>����{�U�Z��W�֧D"�H�w^�8CK�������"��D���<WU���Ko�!�c��
��&jS�o��
��`�Z��r���a��J��8w߰3n���"#Ga����ׁ)�5h�b�o�2�9��Ud�ܱ4_��KEI�1ޙ�x�¡������ӄ�lt&���U6��ܖ���6�5�*ߢ]D��7f�/Y䘗R����"a{9.aT���&w��я�.�/��AJ��ڱ����[T���de���*�p��=��V��G1�??J@/C�	�K12� I��+tu{������S�4� _.��W=�G�W���.+3�A�^ 3�Ԥ��KL�0�K����x<���.�r�=L��'üI~TAPSˣ��e���-��H��d��g����Y$�__O�S(�����eZY�
�����N�(E�<ֈ��݅�hǏZ,DR�co�^�>�&����SV :�\5�ǹ֮��M�e��R:"��c{�x��m���9��#�[��Z���5�LrA��!��Z0Q�hwб��Zqf�����p���k���j�#�B���B�q���2S�M���S���&�GTE���ɭ+j�	`N϶	�ߣ��-NMxU"�@��	�с�L�/"m��<�	J<p�S?^
8��� pY����c�{�u�e�����l�$W�y�A���\-ނhئ�G���k��k�Q�EU�C9;4��SD�P�Y�'r�nQ;!�&���X�m%�����sOF~E���R����>���3f4��������vX��q�����Q�8OE�/��~#��0^ļ��[�~�����j����H��i�׬4��6խ����6ě���,��A3�	w��-�<q� f0��11uޥ!&��(���/��=J1� �X�^<5BR]�`�A隟by?������X0�@��3��OZj�3��Ie�_��;S}F���R|f�鹊�zU7QL��'�Y�����/�t�V�&���S�<��4s���p����p?T����>��g�%Z�5ؗJ`X�4aj����������_���k�������U���?��0���	�r&��o9���۟/��bV+H��h����j�C,�'6�^֙H�P���<��o�S�=�$e�E�J#C��a|3�B�'�?I��"�P�P�|��v��ĝ6Ny��"�F�RY�R�� ����Ls��wŔ���h��vEW��+�(\��Η�oa��j�$F���F'J��^��=���x~:��ۮ1�*�|&�Ծ�o"�W��<�������Ęy���ƞ��|�d� f�"���7�)P&=�ru�R2���e���)3=�A�N��-�^�ɳ��c��aY½���0�T�������%F��B��^�%+�p�C�Fz�(O�+;Di�vey�3	�֥В��V��
0���y�QP,��{~h���;2{��Y�t�K=��e�į��>�~���Ŭ\O��a���#(�L.I��=�У��o��
�޶���l.�"Z����6��u&m��4����*	�z�
��{e���6n����qe�[��NQ��x���U��b�	||Y�>�\�Z��_)909��&�2:�;lu}��pC�a^%�M���n@�Z�����+3E�Nm���|�~!}�R�z��|�5�g�V��s�]��Ҟg'V�U<$F���<����m�-mV��j�6c`l�,F���/�<`[�ԛ��H�`���s�+U;̏����� �ҹe�Ɇ���i]C�B�9D��YI���f
�j��#�-�����)�0?X��Di��Jh�I=T�r��Y�D��&)���Q�#�l�e����)mB���F���'p/ȍ=�#�7��� ���;
�Xvwm�bΠx>ׅ��-���MڼCɈ