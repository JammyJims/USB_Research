XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_>*�;���mM�'���U�P�	)n[��Ԍ�w���H}�6&_!FS����I4 ���
7��Ҧ��(���m��w4OF�R��uT^�sK��*�V��x.������w�'j��o�rX�]W�CD�����{���H�{F"N3?��oC9�z������u\FSa��P��<@U:��	�g�YZ�g�;� W:��_���H���%-qt8�kw�9L�	j6U,���d<W����?�mU �'�DW�[$�NWf�-x�f{�p¯Z3u�~���q��!���Yb�9{��^3��~c��!�oj`Ebne���|p'�"��?6]L���% `��-�6���ܧ0�"z� ��Z���kH��Ƿ�j"�R�Sp-\�㊀����[�Mɋ�M#L����ؿ(��$��%٣?ZH(H>VkӌH��&��x�O��4�ƟQ�k��ۧ#�$5�P��X����&f�Ը,���R&8h��+n���E�K����q✗e��Q�>l���"]�7����0x�3��g$ϯ#0�y��ڷ�0���Z*��	�.��{0+?��9Vٱ�eAi2�pY���/��*S�d������o�^ ��Ɇ}T~@Bx��t�+�#�����)}���P��(�큅���׿T��'-��I4V�����7��Z;�#��"��e�J��BT ����y�r�0������ �H�T�1�$�t�k�D;=C��������E:ڿQ�o��������EjJi�o��;_aXlxVHYEB    2f27     f40fY@�	{�˅�ac�T�rT����*u��#��o�op�s'�S4Fur=J�������Z)7QSȠ�`�o����=�񂿏L����6�`�&m�	�\{*�CPP�B䫶���|��ζ��j'0a8���ܩ�^Ƒ��ؑ�7�gjr9l7��P��!�l5;�FUY�'
^u���3�����x� S)�Zˋ)�󏢥#���
x���[^�!6{04לK&�n?��ۦ����d�I8��`rM=6�ʲ�S�{�yS[�Qc��\�1��6hU� �i17ǧM�X�Ok1J���MzU��3��� z�=���=J�"��В#y�JTϧ�!%�9V�����O6�`(~O���u)J@c��\����m�H�>�:�+����*sf����阻�mü}G���u�}�q{��X47&:E
�q����Oy��.�������d��1�(!bP�9'#.�~	@M`0��'�g� L_J{�j(̓�<ގU�Y쎠TdŸ��x�sO�;���aLn��6�.ʡ��q�8�(Sk��xv�ػ	��z6��n4�	0���%���':+�3l���ȟ�����S��Q�]��g�r���2�B����1c��U&"tL�����)�7�܆�.�nSf{C�
h�Ո00t�lۓ`�6�$,@[��-2f��n���Қr��w�����s)@bcXf����m_q�P/��aw]�k�;4L�Gx�jf���8�cݤ��w�B{yy���2���AK�����@�y�5Ms�p�fFG����S���İO|9 ^@���=�xl���-v�������G_D�#L�.�t�p�=°wB�J͚(>	�MkA� ,�+}L��#�G褰Z�N��>�٩�Yo�C��Xq���l���
G��S�GC�8�V/�e����Û�����J�Ł�-�6���j��w�1g>��		(PU��� ���~0.y�ҿ%���2��>+"��V�l{š@����+EOR)p��}ȗ�>9R�+�^VyӮʲ�H�f]�B�Y�A>7�&��D~{��b��CV6�����,�A"�
ȓ�����-���f�)&��&�&묷�k
z@�<�]"eDzQ�@G�+�)C��ڡcX�$%̀��[���+����}�+5�L��la-"�e�cka�!~l<���N��Sz����z��^F��Q3��� 8rOh���]	��tS�d�m���/P��{��&7V�@3ǮE%b���y{��P�a`u�/ۤ�p %����]q$�~�/�Q36�N�Y9%9h��z��/Q�S�s���z�J�:O�O��!p9)B����j[�VgZeȇ�&�<eY�ڥGPyj���vge�,@�����S~h?T,��N$�h<z�
�
�]�e�o�7Q�Bf�Eaf�T��wa�� :ʼPsŜ�5���Ÿ6k�zg��T��Ou��J��k�B
���'�g4��F�?4��P�^�!FA���y�ȕͭ~$���'��f<$�*=��w�a7���%�;�{��9�G�d��Q/���kIW�8���+'>�2�$ &"�q�zÎ����1�	����iÅ����7>�T?4"�M�G�S� fVfr;5O�"��%���2l*��L��8%|�a+{����h8\pv�Z�-��Gtn�D4���3#1ѻz�@T����O�?67����̴T\ʃY����=��C3��kH���;�|����5 �Y��d���g�C�.�8Z�`.	0A�i���#*��L"�`�kn

�#B�x�I�ge�E�oA�8���T9�PG��W0:�%�/�C�_GIJ�����\�_r�iFQ���������Ћ��w}ٛ���-��gh<�w�3fǞ�Д�r�^ww&�,��m��}���4��L��_��V.о<�lM����%%t{5�x�2�3~��x0��j����1m��W �1�e=!g`���w�L���ۂ�Q��s�y �ߏ�+��)�a(���l�#�*:K�?���+�tR{X�UY �ge�w�m	j񭚒���3!�RgL������0�����"nh~�sG�׉1BF�?��H��[�SJ��CQ*	���ɝvP�=��d���~m���{Ѻ`��7h�5
�@4��m6V+ ��6���YD�x*.ed1;�a�}@���C>b�&�ӿV��\*�ɫ�?���M�֒!�u!Uj��{�����'��|��My��|&E�����I��goQl7,�=�f�D�=���;"�20%(��f���R�%GrAJE������y�d���%��[4����9���?:ӵ}��$�~KaU)g	R�1�0�W��;;$���1'{=����>ug#��s2� r�fb)>����J�ԄmC��)�d<T�"d�(�)��kD6(�F?&��C�4��[8���I���D�]��K<+Ƈ�?�F�}q9�f�͕b�;��In?E��bvߥf�:��g3��WD$\���-]������B]���c�EJ3�Ч$n���i~I�y�!k4~6�v��g*G}'�0�h���ڝ�+-H�F���M�����!���j��ۛȺ����N>�pկ�1i�����O�J �܇?���s��騡I�� ^ ݂��"�Nܭ~����w���ԛ	�nz{�R�j�����$���C�K$�P��v:AQ+�M���@$}<jUw��H�(���ĭ�8:�5:2K�ځ�zp�p�YLnF&Q����"�WK>�v�ʕ d�eQV�U�]�7������6ŕ���#ۦ�i$S�i��
������^)��a9��@Rx/{X��?�胙�Ӫ�
/5oܐx��N>�1�t�Ԛp5o�Wg;�?M.��x�7� ̿������������Ks������m�ú����+8�x׾P1W�њ�g�.Z��?��ߴ�PO�u!�0]c������3#�e�.��_L���qbmj����zA^����@��n���~q϶#(��4b��x���I�0k[�=x<�hx�F:����1�h�Z�ݱ���a�˂��Oo�*}&,�^�������@e;��=r���c��8L[��Q���4�1Z�4���K��+���P�y�ޥk�⿃V��%��$�IT�����|�HI�e��*��T\��	i�k�DmSl3%��-�⇑��VU~ՁL<�z��n�"k>}�?�n�/�Z��!��k(�D=�X���\�S���4��52fu���៝�I�Ѩ�cٟB2~�o��\��5�	�b��ŀ�����q>iӱ	5�ӁqF	z�٩V�`�򰕫4�3]��`�?~�)��>�PJꠍ B���`.�8��Gzx��c�:�H�
`(�`���
=�ٳ���=���If�I7�6�*OpS�ԁr]�6D��/k��|�������F��c��Xh���\�G�`4Q�oч_硥��������r'���!h�����f~��\�J��y�����-����&w0KH#T�����6���� g�F��˕P?��?VU�z;�i��s�t����]�AbT8k�Ǡ~$�>T��JD'.a$��Lج�&�@��},x�˽��[H񮠑U���e���̵�����>�EQu�hL��r��C�Ԫ&�B�0���_����|s�t���f�����^��;�6�'�$���F/�B������*u�fĤ�qw�g��6��b������$��0+4� iWg
���i�����H�a_]V~	CŉT�5����������Y� +�QO�4X�1�p?	0N��V�P�C��'#s���,�ݞ1J�U%a�×6�s�18�4谧�"�]�'���v&�)i�C��6�Q�a,^A