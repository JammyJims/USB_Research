XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ZNhZۜ<<�De%I4L�[�O�n�3 AM��7��[�&���Y�}������~�t��n�[�-���v��*_��lo �ðP����q����1+A̂9}gTc��9����;N��Df���\za`����E��|��SX��7���,�����]`����M�פ�Oh;�Nl�$��3Χͣ�f�9���q�$-�=�d���l`�����18�B��� �c|$�oc(r��yNU���2N�CR�H"2Ь�W���|VC���y5$$MTT&l� �j�+��~�@�)@��::��5}ur'/��O��~��u7�T ȑHF����f�;���ʲ	��UXP`�\��ɀ"\g��h��ĠI<}���HS��8oz�O�ը^z��2�ż�����d>�\��������q�-�3����E\TZ�����3_���Ɓ�I�؃���>��R�[�/2���	�9����� o�O���35���l;��|�\��}������d�(�t�MԄ'���߃*���[��`,�ɑ��R�s�%�FI	�'��N������F�?�`���č�h������+�Q"��{�؏T4v�W�3@��}V�eq��@0���#����Xc|��3x�5��Q�y|샧F���AhN�p��K����h�
Q��F5g���L���9��ƛ�q��x9�3���R�e�btQM�s��9�.�)ϒ�=}}��JE)�%�"�XlxVHYEB    68e5    10b0(Q�v=[�o �5(�@�m{X6PNX�W	U-�� ��@u6�՚>`:~�[�ŧކt6]�`:�	n�	'�d�ixMڄ�[�6��ުR��{w���;�-�H
�R#���݅m�⎩����8��������mc�R�f�8�v]+�o~Wm�����<N�)��U#�Ii%��; ��UB��9*�ؘ�y	�F���[D&Q�bf*E^eN����謠��3�o�˦M.sC�t�W�e��,ڷ$i�P���c*�s@p秋���^�q���7Q�T~��G��.i��^Ӊ	.G�4���T�F��ȋ������_�h$s�L��i#,�
��5˯�W��.�wR��`�/¦�y�C���Gd�7r�[��~��7�2��d������K8g���1�=�6U�����ܧ��'F��$�:�E���f�m���3�c����||m2(�-���fRn��ğ�����Z�u!��2�-���Q]�:`�}�������/����'��Ӿ}y�z�u���߈�P�N���#�2�A����/����ҏ�~S�n��S���,���	�>g���[ vd`��P��U��)��f�9�YmF��qxE0�?�ۆ��[S۲����?�dۄ<�5S-��E�n�!�"F#�e�fϮ�-V�	��;�F����P{��|tx��ʌ����|����L����[RD����4H��V)6�R���`_�t�����o~<��Y�^H�3�O�߽��J@�����{��|�
\�$���iʶe04�h5,����ĳ��v*�+��%ǁo�KfU>��"���� 8��R�=u2,�����K��c�~��������$�4�e��35��Rā���%z�3�3v#�6�D���Z� oOFu�8�{[��2�I#���Ѻ8�T)^�N�An:���#o��H+C%�L/.�c���iRT��)z��e=�T+�@e��D%+u57[��-�ٳ=��t�2�-1�a�lV��-%������\�0�E�A�ᓈ��B������,�����Ʋ~3<|�T�P��v����tq����N�/��U-e�ٝ�F����@W����R|������8�͚'����¸�q��4�B�~�9��"��H�� P��t;�Y�	:��n���oldZ���3�����
�����L�5�R��V�=���<�g��u��;Y�~>I�%���� ?�}���T4/b{�?ӏ�OJ��x�t-��G_W��X��o�p�'o����j������f<W��[�2}�|���@��Z��р���!:X���5,��@���F}�C)%Wʮ	}�G�&PE��luI�Į,��>��z�鼻���[�W�N����Qt��_,�@�{�z��B��0��˽w�F|��� ;�"�2yQ �2�%h���WY �r���5˚�jxE'>�k�pu��Y	b��hN���i����s�3c��(�yd�(&�U���'L7l*4H8�ע4ԇ�w) ��~��t���v�E�ȣb^S�B�������\³�1,q(ZĀ�py����q��,�?�&<�-�w���u�$Ƹ��Kΐq-�㗻w��2�Z�N�A�ڱb�C;C�[ﮒd�����G$V�Ǟ赗�h;�b8�J�T�!��	�{>�Qx�0�_��A ��x�"��@ ��{W����yq�G9����1�N*����/�z��d�b(̅EfR��+��A��T���3נP��ۨS�o<���L6Λܦ��H����i�6�[jE�P�:�9|[�ǪB��ӕ��D�y}�	��)�K��֬s�l�%����%�6��F�������T/�@���Hm���Tfn������/C�?��+}��WN��ѕ�F��4�"e[Ļ��1�%�<��_	H���C H���7�����+~�j'v��/�ke9���������E^Z��8����\z�|r8�0��o��������K�i��[Gv�({�ۅ�,%��M�R@�v�yyD�"�|.ߟ���m����k[�E��,�J俾^����:��_ŧ()&NNR5��H�Q$&���{H����x��j��)���ajX�\�F4�Fv0x����y��� y=R���,v��_�v���\O��p����r� �o|;��\?���mvD�[�+~�X@��e&z;IF)�sȻ۳Ե�fq�Y�w>�b�۸�0'P�o����zS���#�,4$7��|�%)q��s�$˕�cۚQ���s�����R'/��f��ly�S��cz�"��gS���_%Ҏ��K�/�������k;^a���3l�����U=��D��2nQci��HM�!_��}j��np�E �UXu�����_��2�9�ɹ47�$wV�P�r�l����W��x�?ޢ���#hA;'�;-k�>g66�8x'p��2�$���.�|�	ry<������g�-�"Cz�+3���t~��K[�w�L����o�7�	�kD�[���EK���ﮠ�}��Z��	\֎*�����������r�y���70���D��R��gO3���._��q�QL��5H��I2~z)�=�ZMOq�#(��ݐ�3H�3>��Wj?��&;H�w�4C�s���@�t99$չ���X~[�YK����+�����ٍ�E!4oSù���U-��s�ܞ!��h�=�~��*P�h�?�&����h&��ND����j�T�h�� �B�i���.�>����s�s�P�L+e��C�����5Eo$��>��@Жys��*����;�F-���u��/!d��	�Զ�z5.��i�Iiv����"���Oٻ�t��wp�*��nmC��� +�+���z�iF�r`ܟwZH�.�����W1:5t9�^Gl
�5�����%��n58m{��l!Í{L�t����38���.��Uh>-���Ū.z�0��p��O��HI�B�����
ɳ/��������M�����\�х����q��Κ%�o�ۤO�ϵ��n��M
�gl��wv�����Cq4?�Ks�s��8+�FRʉ�Q���Xa���_o��Z�xe�/�R��*�Y!�>ڣ��1>J����=��{� *Y�Mjd3
���& � j`�B�5n��0=��,�E������rt��τ>�o�r���-���K���{k��K��b�t{obvA@�u�d6d��1,���a�r��'�o6�fH�+��2�" \��=`��m��m ������}�SY_}�e����b�<�`ˍ /y�y��+���� "��Ȟ����jx���+�ˍ��( H����9&��Z�RfO`vCቔh,�Ȥu��ԃ�_�P�x�޽��� ��p�4��#�.m̈o0�v��`�U�L���؟m �#�öR��S��N�����en�bku���Kb��D�#�_���K0n�4
@�B �2z�r��y�2v��x$��4$�G�%O�b�'�Z.����dL��а�H g��?:�v)�]��֞n�j{�FS#ন����2 �_���.#�;��0C��(���d�n+�qW�w*�A��.��,x7P+M���U7R+���a�mԳ���7��>����ے�i�=�$/5��7J����G��SUH9�K�ᐡ׹���BVFO�ŭH��7_�}F#�x䢑�8W�V A,N^�B�H���#k?��UA�B�i[�;��(c��	����q�'�Ǥ��x1vU�?��T�ʳ��N������}�^���ڷ�@Ā����gcS�iP�x9^&E#����IE�2nB�kU���>8���zW�,���{#����-�D	��Έ� S�'�3eQq�¶�95N����k��1�nv��� ��_�J���{��@S�1��E�Xe��ԋvq�$�Q���"�Pz�kH�����Bg�3�*�D��'��E������o��C{��t~��#R�XӒ��:!	���5�l̞SWe>�����Ui��ށQgWy6�n����T&Jf���]��hb�)Ƈw�J�g}����d�09���C�E|��!1����-�qs'ũ��!(E�\�r�P�M�u�NZvE���p���;�c��{:�=���YAFe��k{x6����q~zL�i�zKjjx�Q��