XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z>>ϳ;\]���䧮ʢ��R����fWw=35#V�H��O����~Awpb�ևW; %\�QP	RA�1�l����� ���������w�P,�~�|�g�� 977�t�թ$�j:uk�pYÌ#n�<� _���@�,&�:��!��=���+��=�z-N�Y�Y�˝�([vh����7o�{��ϭ�� ��.z���@=H���?�:�U�(���Ho�H��&n������!�v�P��g���L�0�.,���R�8d��l�9nD���ys��_���!Z�����ҕ������p֤��"�M�p*���-~�3���C�����m~|���^�xG��(�X�|�9��f� �A7��=�U�@�W�q�5M�$�ݻ{X��҉����������׭�,��%�X�7�8��z3t�~�^�\�����Ǎ��ḙ��(��2!��ܟ^BQ�V��2ͼ'���)��:���"w,�`�������5FAA,�j�x�����/�a��v0`�wάs:L,ևCϬ*3��p���R�~h
`K�Č#�Ҩ|?�� }.���K�J/{i�h��,�����nVWw�'�V1���J��[��g~독 ��]JC�ɑ,�@rX�ڕ�>�!d��FrX=�?�pl���t���,=�Z�����d>��Gr���o�!<�D�W(����[M��o�:�𗳱��ณAX����Zÿ�y&�e�����/�P�#{�&(�XlxVHYEB    463d    12e0�$Y�lT}��N܁�u��� ����kt��������%��)-��k7P�j�(�s97"Z]����<(�9�O��d+g������@7gd&�{�����Jv���8�0������m��d��V`r����*u�w��HIp �`�ul�Y����J��}�<a�EvW6Q����Q���{�|^�@���-2��c�S	R��cv�0J�IOV��`��H?�磷�Q�677pt_mEh+������#�&���������2�E�C`�[�ms�Y� F���
I,ip��0�A<"�q�)���v�'��Y�Q�.d.Eb�Q'6�aѷf�a/��H���k#�)g�����W:f����UxT<f�
��@��tfN7�j~v)r7��3;�j�Sٍڦq��m:�w �����@��s�	���b�H���B_���[Qi�:�W(Ӝ���E(��'�:F�������|�-��1^�RX��`r�n�|���P�G��sU���`�(@�h����B�G��8S���5D]�υ�X������6Y�\�*�2�(��s��a�\�����y�ij+�۩�����X���X�"��o���,�Oꢅ���oJC�,B�9[�K�6r��V~)!3������QaJe|�G�.t�"�4�M/���3�e�}�s\^��4�"J�/�����\X�R?�~�$��t����m\�(�S}�Ni��3	P/�s�p���6��'�*Ciԑ�k;:�VX]�]�G��`�}U��q#5^�̭��Ƽȴ��}��]3�,�������˷�#�+RS�Vo �:0��Ib�oc��Q��^�?/	�w��Y�VKDŰ��E���q��_O�6E$	����(���^&�?ΜP�D�ϋ�J>�˺!�L:$�v�����YV��4T�c8xpx����D�eF����:mB�r��M��l��]yS�$O4�g�]���:���*��Pv��=�B�������Q��c
�%�d�,���)�S�(|X�J�yNV��]��꾰mJ��p�ᡗ���,�^�c
P��.7��4'6e'��9��'VO�b �?������������ds���0�nH���/FH�
]�(0��8�C����(:�N'?����[���pe[
��Q �u$��i�����@ۯTJ'� ���b�������ϼ:DDr�t����.�
�C��~��$�ǵ��ݑļ������A�a�>�O��[G~���d���~C��ly
YU���?�$��P%oz�7R�~�cH�Qb:7(6�Q�M�d��Qe�Qo&����D?�s��Y��c�8؝|0]i<�R�don=6(�;��F�=gz$��?�k��!�K1��d:Kou� ZE�D9)5��V���}�>U[�{��I����&6�=6��?m[������|�PcspfG�x��Au�]�k#�am�)�1K�`���`S�|��'#��X$�P��yԉ�{�xV���!��O��:��pݽ��y�IA�u2h>��K+���Nt$ �2\�4�+�B��HǏ����!�E�bOW�sڬ�dT�ǳ�/��,4���<rH��V)e���YR��js=�vI���0�~fS��X_ζ!t��k@^Kh�q���{�%�b����б�7ڷ�ɿ���+p�uSV���$�v1դ��4W����X(DIf��I�G ������{�m3� �����wĮ�|u��b˙6S����ʾ�9���7�o�Ef�|<�u��G���S��?ο��ڹ��w��mhhlv�
A��8�#��~��ĝ�^u�>嵴&��������W(PH�Y��dlz�0�W%�5p��I���T�XH�� �>�k�M�ۍ�����X���`���o�M}Ɣ�7]sU��y�%���0�x�����u@�My�/�������OÌ�-�����Ue��/���ǽ�*Y+��J��kj\͆�Z��	�C�<i����Z�����5ߙ*��?�b���=�QΝX�Y[������Fβ-��0�c/�³���k�)j�@�6�YإQ�E���������fBEc�k�ޔ7�n3�������_���2�ё�!F���:%3�� ����v��|�F�i�Y&��xPNL���O��ˉ�6nj��p�4]�?ZH:�r��z�h(Ϻ�	sX@��߻ʩO��^�Lշ����x{(����â�a��lh�jk��į���H^~t/is��x�ww)����dr֏�!��?��RĦ0�{�B�$�lw���a���7j��AE�n�S[�JZ��9{�		���O����Ʃ��J��v#�#��hi�y˅�|���:�U�ڴq�����)�2w����4�v���a;Z�;!C�Iq��k>�uV?Z�^���ZSW�\���v�fo,r^�OM�,κ��wT�ڏxXPN���%[��l��56��p�T%Rë��R1��W���􎴞�,�H����+Γ�1�	/�ͩN���C��D�W^*�B��Mrd��P"��H�V�	fdd�e��)��Di��r*��%��Dç�D��}���`uK ?�I�{.0޾E,Yq�����&ݐMe�S=�ơ�+�ﰍ^l�]����U�79ijǐ��WZH�Q�WnF�^u����6d/�{�d�du�f�>�AL���&7g8�)mv��=����wk�k���F��:م���N5�^���JD�(ZV�.�,4i�e�C`M��@]������$2��Q���ѣ��VГ��X}6�m�/K�[��57j{v�a��^�o�b���W�(�Mˁɓ�NK����l,ޘ�)�;�	Mjpk�㲢��|��C�$~i����΍/������s�&�.O�Qx�оc�V���h�&�A���&�-�Dv��J:֋q#��|����(�d�dw%�	p8�H�PҪ�W�mfD�ftX���$��@��p�-@�+niz�u���#�!V]f�RD$�BT�}V�=Xֵ�QZ�}���w ��lR)ȗ��L�hlM:�k��E/���N��5y˓�RԬ�̱-N'��׺4b��D(��&����2���L�b3H
��;c����>�*B���j�32|K��}PH�&�n5�&�4%�$u4��tr��!%��1�@=H�4�:op�^WR0��.]🖾u#Q��d�3
��<���� <��;w�U.�a��K��oGq<�}J�')���t��ge�O�L&�pp3P�JK��R*�Au��_m��N$�����؁h�0������Q��V2ü�4���s��pvjּ��iU�����,ۂS�R
� a�/�hʵAB�6�r��I��Vt��
,P"�+9��`>���M�4�+��%�hѹd�c�&gh��M�TI��k�Fڟh^z�e��u�f'����˯�P�Cj��܊���1 \	.�A��|O�N��d�{�����Ϧ�����<%�3�Șq�.$M4��y�k����Df��:B[r,��c��Hr�M�0�QM��1a2�it:���"'X�k��B�|8��#���7/���4����x�p4���J�=�Z���n��m�]�j^�}����Z�)�3��L��]��?����r�8��%�
R��M.'A�2�Z������d��F\�yV�05���Һ�����pT��p>����*|��4F��S��`(�V<Ӕ�B�)���@qB�/�$��[P˙g�}$Pm|���?�b�������0�?̶��E��l�<t6�p��T����8����j7W�ݙh��2�ؑ�ĵ�]GX����H$D1V��޺H��,:��#��*�ȴn᜸����m�	��=��P[BM%c��R�V6l�d̷R3��������˪�|C��/!�JJUnM���i�.����v�aqͻ}H�ckB��謒�]���{�C��(/u�Z"�T�$5j����fP��3h���*v��}�媉�_�u��{�-��I[�Y������D�p'��[qsՃ霘+/.iR�i?NI�<��S�`7b�qn�߬BZ�Ecs�L}�r:��IP��Z���w&�c��O�y�2�"WH8��s��WN�#?ǀf^�� @
|��˽�����Q7Ɛ�J?�f$��ǚ}���n'��|�S	8k f��:�Ǟ���p���c�N'�������v$�	��p%$����sEt:����Dŵ/��-�(s��`�H���C��tS��Oz3)sƲU��nL���KD�@�W5�wU��PF�dx�w���u1����:�%�O�K�t�{�����u�8ʹz$�ܮ�cG��_�O�"�$�K���!d>��,YQ�)O�^ҧ�@��[���nx���
WT[Z��c�V�|��ڵ3������,�a8��2���c'��G��0�dj�·�:��v��W���g~M���Si�&�-��V�:��g�ɥ�(h�nK�0S-�Xi܏�Yt8��}%�U�n�T.�-�N���8�#�[���5��p�2�}�FA��.^���<���ː0)��T��FG5�V�{^���D����Yy�_E$s� ��lz�CVȡ;e��Y1�(��Nr
�K��@�f�МcH��*��42°��s��Y!��LF4�R���2R��﷮�6�5�u�60�Ō[G��m
��q(~�ro���f4��=Z!�Οe/ys�a�܅i��"aPzz��}��#�w�?��;1�m���cM/��v�X��T�%z+צ�N�W�*l,�p5l?��y�R�Ww��iXҐ.����n