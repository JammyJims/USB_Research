XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ЯǭD�">{�����؁i��V&�'�^���^%�b2a H��p����U��A�״bt�}.3��
h6���G[�kj@��W���-i�!�E�k���@�e�gbJ�^�v+9������@�*�KDzx?$!��� ��Q�d��cS��R���r!�z}p�vTxT�gȏ_ũ��=����B�ڴ+*MW�ʓY��u�fI�>�J�fl�TK���q�/z��s݁�r�������M���d"7�'[6Y܉�VA�Vt��W���y�j������@-M2�`�j�7�F�M�h�|��d1��Ӭ/Un��1*4��;#��݊��o�E�?��-�x����^��'�>�S�E
�DI��0S*���lBk��0̀�U�'+L8��n��R�!����R�0e:5(Y�3�K����*T6k<����1����H~���E�xX1|�b���J�'�d�	G�eZ%2J(�Xu�J��3-��xo�ʈ��L�2��	ɽ�4���Pj�b�����C덑�Y'���E�Z���K�{���X#��L�0/R����ˊ�I���A�Ú���Q�#*�������PŤk�7�ayd�Zhm(����������,[F*m��K|�7�Q��'�v�7�+�E��Gˀ�y����Я;'��/�����y�┇͒>y�O�=s�
v�����@C}璾�L��tg|Z�1!|Z������f,�wzj݄H��]�h2r;pN�e1�'� A��&�j7ge��(�;XlxVHYEB     97f     290�{�{D7CX��Ru�D!@���[�v�B�����{�WĔ��J/@�x��p��"[6��\�
]v�$�q�k���fĕ�y�^u��Pb�ۺM���v��R͵�~FR����*2��q�`���Yb!���)���D �'f�����T�?��l�V���8S�*쩦Փ8�4��G~zѥ���M�F��f�`�|8���)�z��S�`O踦��}x��x���%W�&�י�Z�{��k��g�:�b�%αޒ�2�S��.V�: w�w�0DE���ɱ�Ŝ K��'�)*SX�*�SoG"��w��}5���$��oHkeJ�qH��~����b�i�[^EM��/��OӬ�I����"�:�C�VGO]��� ��3:ݬ@���|���$�dv�>���»?%0���+�W(��3���v,t߀���r���L/�G���S���F���
��"f!��Fq��%�߾�?� T� �{�E�[`�vNd���`�8ԗ���J�-�٢��Dl��}���uG{�XJ�@E�mx%$�(�����R���n�χ��£��鸺�>�A�^@ӼQ�"��Р�OK�;Y�[�G�	>�O)�j��ߚ2h�M���e>&&D/�Ӿ�/`�mB�i/