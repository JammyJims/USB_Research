XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j0#_|��nu��V{�o�}��Oj�x9��i�m� E����`,��u �J��܏ [9�XfR��^W�����3(�jePT>r�t)�K�K��[f]��Of��
�ƀ�Z,������H��Z �� q�6������p�/R�ad��+���zR��~Y\_��9C�-�?>�}��<*y�<h���ʖ���1����b!�,+J,)aJ9�EW++�[O\̡X����L�v�t��ڠ({U��9�Zg`}xt�a&��g��<�`��������P2�m�nA+h1wT_��{ੇ${8���(0PƩ6��F$�/@
A�=��(F�C���4�c��Q��G��^���kH����*�,��=��&��'�k������a֔��.�M_�_V<J�Ih$H��L~���č����a�x��h�~���_��7P�|,�Y_����b�C��uO��X>$-��B>���(d�Zy��g�	I��,�Z�Δw�:T�����;���$j:^� LO��"�~��~?��Y_�8]�M������2�N*���)����@��sߏ�)g�]|w�F��|����]�~����X�_����0ݿ��,Y��]S��̷��,)��8���KxW�� �oD���@q^�ֈ bw��{�T�r7D���S��A1o�����:8@M�7r;��*�ʆؙ�]���X�n��59�ѩ�_��D��ag
�e1��w�4m���P"���|]��mf�U�h��XlxVHYEB    18c0     8b0!������i�Ghlx�V [f�7o���O�I��!0̔O����z�𣋻�'3��h�i���Iצ��@i�"����xf��Y����!��Ռ�\k�d�>��:ʃ*&� s��P�����z��)�n��.���#J�>W?��o:�Fw�����F�S5� �X[d���sVn�?L�<_t�����~��e��<A�v-b��%:Y��;����}wb���͵L:��j�B��s�3��݃���2��O@�1�S�J�fA�R�W�s_�ԝ�xX~D�fi�cuF���V�ކ8�U��6|�p��&<@%�����݋�;�3�5=���:����מ�́_���:���z��T(,�ð	`-up���4[[ud����rl��ګ :�Rj��(!�X�:���,�y���m�-T��f��F�<#��Պ�ꄕ2��؈�Խ��[dN�}�i#���qh��m�t�����>^�bS�K�	�كj�k��!;��#XM$o�[�	BS�Vw;5���T,6�A�}�{�Ex��F�z�x-�!������ �`X��kY-�곦ʗ�A�^�J�����|b�g�Զ!��@��s��jYA[���Y�y�n�K�)��WŢq-W��c�\���6t8�����0<D����<n'����h�.��t��P��í��"���]�c���x�L���7�;��ҝ� Gz���%0.�b����	ke��i�|��.��1W�����H�-������al# ^�4�rp��;����׌x-Q��R�+�(��J���K��5	��2&9�kr��ɕ��J�Ts�w�I7��TaGmlk^i*
���_��	t���{�+1,�W�͍G�I���Qv6�q_�g�f�Gi�"�6Ǹ��������JL^�5���)�E$�:���hE�Ք�{V�>���[N(�K��ƌOd�~� ��ӣA���$�k�=��� 0�@^�І!�^���\a�Xk�+��U�!�o�ݯ�R��$�����lߢ�ȑŁ�H��$H�e�[+��:8
�
��l�w1�5AU2����c�\�J���K/����|��/��ۿ�f�3�yV���T%IO�Su��w�\,�e�����, �e����$���Կ�'T���ȟږf�eYOV�e�� �|��Ĥ��	Zr���,4�M����>�_���q�Rq�k\
���B�|�b���w*�CF7�8�lbW���r
 E��c�^�w#�Q��$�c%�(��P����
6�Y=��u���^"�lE[���,�\�౽��<��c�y�g��=�x�d�������$�(�e��GwN�==�ȎK��lt3�x�DB�����Tm����djz��]o�k|<G��[��)����/�܊����Ⓦ�G��ܭ�&�a������e���Z�Rs"�hj� M��&��6dr+��gQ�rֈ�9~��[��t[������|�&�O��H�rt:�S��:�W���%�O���$�#������:~{���-ʛ�H6�>"�����M���Y͕!�:Çh$ձ�dXn7�	�
A!]�׾��+�,P�c
�J���Q?yKP����'�Y[F�K�3̐F^<u�_�KG��Ѵ�~=c��6|��S<�Į�K�T�����:uL�Γ���Xy�������R@�Ƿ���P*�x�	�J[K���K+�b�(7���a}�=�/�������@��-F�s�'�yx��J�>;Q0K�9�����`�M��#v�_��&ʫ "�Ђ��S%���ZT����\��i�_�� �@:]����nŖ!ׁ��}j�r�����-�Pq5�Y_�L3F(���
�ܝ�0 �K��7%�z4G�Pڨ���wɮ��hx�St�V����ms�x\eV��#�w�,;ן	(#�~	�#�l��9�m��郡$P��B��_I
��TM��$��7�cy�R�۠�9~'��Zcd��_�#Y6�m|��rr���4���⭗�mq��k�-�����ǘ �]�$����MZ�8�Z�+E�s�$�@#�ϝjg	nG�Aս�X�A�&��;�5���s*�h�%��@�=z����w �ݰ4���s�k�B��*r�#��3��}Kq����ĒA35��G��sZVa�і����o:V�