XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v���v��F��I���?����}x� z�!�Xg���*��;�����&�v�7c`Y�h�n�N|������|>�)�H�JUܑ�8:�H�iQ}�2�G'��L=��}�Y��a��K�<0��\���Ycu�L^��e-q&�E��77��Y�E�U�AB�]�O1r��\�,�(�᝸_��7[���I���;�3���*e�c���pBe����Òꍟ�x�-G�Ɛ�d,�����,⯼��(|��������%��5@m6�D�"&��Љ�BXOV��q�>4���7��&�JS�t�����qIOM�C_P2-s$I��Ų�y���~mwX����`���gd�
���%��͕��lⷾz!�GIϖ�p��[K��6�F����?�9o`�;�@̓5�ɳ����%$?�>	�]����M����2�ҬD��a�����n)�����6�Dyۍ��`�]Ǔe���$$ϻE�,�����i�X�0�`b�����d��JP�q��4Y3��v�k?�bgu80�l7)��q�_�_�);6�2����}1N���@��_k�qx�EϾ<���pa�.���_�O��Ve�j�jsd�U��4�:��r! � ����g�� "�Y$`�TZ�
H-���0��G��[X�m0�hF���uep��E|4��t�fK��R3$�	fŬ�/" *nx���`��{o�a.9�s9��چ�-��r��JO�_�׸a��XlxVHYEB    9ef1    1a70��wu�{JVN۽�V������i�
.򺗄�$�a�za��a3ɟ�9�!�E߽{�&���,yi)ߓy�����2}��r���}�.�%�.�r��SXM�Q�>���a���ۄ�=؏6�x�x;��3��^�E�g�)�4v�:~Θu~C��5[�?���؋���/!�h��� �_�}�7V ��Ή &����Ci��'}���J�.�����$&�D@Y|8]_�H��*X=�b����h������L�������>�Q�Ȃ�!���:�&��>���D!i���~ic�XjFٻ�J�_���W�_��̈́�������(�C�Ɂ_b��L�uˆ騷�EH���C/�uhv&@����2-����MOF� -8�
#�T�ca�[7V)��a���W� �|`�^=iK����r���֡!m1%}��[���ޱ� �U��<V��D���l&���8��<�-<A����=��Z���i��T�!7��t�F�Vq��-�H��`È}Ye��$����X3���u��շ)$�RI�o�1_X��ӂ����K9P���w<Q�s�ٴ3��d�`>���3�ˎw�;��͋��7��P�2�V5�n�	[����J���E��4���U���}F��$`����er��i�G1�y+�6{�q�$��h��W�	�Q�QM+�5�g�"�5�O�;G3	z�{r���]P�**���(�`1D��%�u��5�x��A�G��SuM�V&�X�$j��쒟p��hٸ��(����𭀓��"�5w�W3~��	����]8X̫�A>u����̈�B�9iUB�z/�jn��G�M.�I����z~�aBln����ԥ��B!0���R�	sQe��R�������7SC�g,LXUK�%���^��j|��Xo��Df��w��i, ^t����ܴ�Eew��_��y&���~�j ����"������<�&;����y�,�~��<+�<8hm釐�-2��Q�B�DC�\���I�t��w��7۶��vm��YI�E�S�0Wu.��Q���c�#���m3�f�l�V>c�LT)��n�W�Ł��	/��(w���#�!���"�t���>�W��L�x��r��Y��B�}./���7eW)�b�}�MT��[W$�G�Ͱp��>]�Q���$���m���fϹ.�o��0�``�&�� Q:�05�ߞ��t�K�tī�s�:㕽6��E�d
 }��?���������n����k�����&�y�F�Ĩ,M;F�k�"��E�o@��c���O�����ʙ(�O '�VJ����CwO�ΌKU�p&j�W~<t<�؀��O�x;1Z��谘��W/
���#��by��o�p��x���l�n�af�=?����2щ��WnDGHd�fyv�&���v��� ��ZD���^�	2��s�v�;��U���/�?��=���wp����h��G�fn������# �Vz�!���~�#m=<шH�;�������Z��!M��%ȱiT@.�Y��Dֵ�9�s�r��/��I]��'�^]�X�7	 I�-�Mwӡ(b�I�c���H��$>� s�ɾi�C�jwQj�{��z8c��%�W�����Eu�-uc:=������g��L�Nm5%�N<�w{(�C��)ϕ���wh�\1�@�q��
�u��(����P���诔z<�K�����(��Q�/ �ފ���x:׸`�}�:�wDypU�z�T�a��W���7)~A�̡c����v���6^�t�&}\�g���=��%*h �߅��x�hxG�!�$6*�j�rܹ0;�9��`H��/�E"hHC4 ���>u����}sX�`��4H,���s){��b��'@�6P��*���M�!��J�����|>�؀ƥI󰗡����#4zL_��n����;�}�D�咹pVΙ,	�C4;گ�{�ū
]q�϶���:�'�XXRA-=2�	~���ڒ���"����L4(ȸ�	�-�7xe�s1>aTY=;� no�\]h���>G�7�jzP��.��(Q��D�$�V�O++5"��>}NئV(���Cy���aD�Ԗ��o�o7n�gD-lf�������:�I(��	�쐵̻�A�EZ�� ���\����*��w7���s.L�ziS��ѮDR�<dK	��a���/W!ˍj��dyj)��k�x%rWٚzP�X��_i2g[S���U=FK8/�uv��m���_j ��Yj��l�P�Ya|j��DG)E[ �Zc��`�칝]}�I(�I7`��Э����&��"Ʊ�1e�[� 碏P�GΗ	����Y6�d|�H���H���u��>��(����ջkJK�r�Ū8���
j��H�l�S����{p�܅�m��	/���?ĩXW�d���t���/H@\_�,�큘��'�H�Z���.��8��3���a�� �bS�p��lN�f?��$�]��@�S�J�eT��A~�Y[�&g�'E	f�����y��ֱ��N�Ă�X@Q���g䇘l[��;(�i�-��1��j��V?���'��v��>z��]		眶zC���:'���bK d�b&�DT=9�~�E����|���A�f����@t������Y�2u	�q�W̧ ��G�Yo,��|@���WO	���Y��|��c:�U;O{���N�2K7��0�uԸ�]C�@��?��BlP�^����EG޽��K�,m��V�x?(+g�]��o��ˁ�kˍI^;���WtK�&� � �E$`�U�����b����^Λ��ڊ��,{To^��W�D�
U��W"��?UώU���6F�v�����1,n���5#C�YWV�+�	8����@o�Lo���r?3��UJd	�p.�h&���w��q�Y �(�������)�;䨳�'�1���l�3�-�/�c�o�Ѻ%g�ozXD��"�E^E���3Q��x�"c�O�f{b�.�������̬��W������N^f�D]��5���0$@�'�[%d��E����'����;:x�İ08.$ ������T����z��A�E(��Gk?�/�uv0~�9h���]���!�<�"?&��yc6e{�bSU�� �t�H��Snw�%a���͝k|���F EYK3x�Б����5�g����0���%�-��7�ٌ.�v!���RlS��� s�O��X����������i$���~���:m�
��l!�)�
�V�u��� �|6X�j��>0���Z��I�{P�\�9��ϰ�3lޘ;e
�Iҫ������#'��_��/��X�̓�a�Tbj7&�Ȧ�_����p[����'��L�Ҭ�"3�\H��{Ό��w1&U�&��K�޺��k�Q��e�CꑐPZ"-���c��u�˵B$���f��|�,�r� ����Y\:�}*�,Mg��#�{L�[����[A�����9�W���� �ԁ8pw�ص0�Ow��Vh��4��q��^O�[(r ���^V���&e:���/8J�pF��lگ����4U	�#Z-����B́�	U|�/�g�o+�b�( � @1��\S�D��
��?	�����k�,q�'�Iqʲ/�b�(�����G6�l�'�jAlo�C���3���7��lg�� �Q ��]���Ed���SKf(h����!����<�N�Vk�oo��.^" 
�k�}�ӹ�抖�-��X:����#ռ��4yH`,��On��>N���n�"P�E�����A��8:9(��	*=��M��W��	bd��p� 8]���^��.��I�ѐ����y���P`�P��M���7�"�Q@�̢�מ�=��Ն�]_U�5�Qھ�/|��A%e<{&�aBR�I�J��1q6[�M)`���e����t����r q�����{R����i!����h:��{�S
�����K=�UJ���$ϣɾ��C�	\����iH�T��އ}8������*cN2	2��Q�����HSI� w���X4�{)��H;��[�]��#����Y��ɠ!��f߲�*�%��L�sƆ��>�Fd�i##?zFhK�GP9�LT�'�n��2�KC�=� �A���>?B wܯL{T���*�م`{��scy���S��B
�˯:u~�⤐��=���x���n�w|��8��R���,Yʎ�����?+!�/I�;����<E�[�*qa�A��n�c���8[��ǽ�q�� Q�,�f+-����, ��8ߓ=둷'ԃcVy��g��U�PH,~t�H�ӷ�'�5�b�=����E��\?ޔP/r�ղr��Q�j��V�}�����3��4����>v0���Z����zm'���B#���e9��(�	

��7?�����I�
�V������J�����x:��ۆ褐6#�oޱ6m�]y���O8��e��Ue�6t�I�Ѕ��^���=k&��v������.�Cs��߃��1	Ex`Wuƒ�v�Z�$�AE���:��Wi�v(�^�a2X����a"q��R7֏�]����W�^ ���0W��~y���.V ~��S�������vZ��9dD������p'p���9)o��C��ܜ�i2��D�F\������������8��:pٹO��=��j-�\������Y��A�~:M�6{4�6��o�J��A��+��\Y�!�g���̢�o��ݡ�вE���Hٳ/�A�8W�+a`F��Bq\�	�g/h�wF�sr�HV��4X��v���bDG.
�Y ,�L��U�Y��\// \S�M?�n�R6C�&B�5!� �.Ig*�?�MTL��,��\�������2�|���2����l� �Q)N����	
DJ�!�.2�(i$Ոh'd��d���;,�Sy�����`I���bȣ�[�\����z�Nk.?��7D� ����dAQ���"mB�>8�.9<GIh�j�Տuj�h���%EH�1{�f}��e?k��Һ.�o8[֬p�o�ʩ��T�f���{F�QW��ӯG<���ۏ4�ݠ^��*`3}Y,�>�'�	+��_�ǩ�L�pD'@a/-�8����?��s�E
ޤ?ׄM|�����	x�Q��Ǿ.f�#"�Xv.Ӏ�x�fyr}�j�~�M��+�=�v�^�d�^��}	z�)�8�g�2Ya�s�#�%g�핀Ղ������y�+K�D�}����+��ꨎ:���BJf�P�z��`
�j���V��T��/����.2F<��"z�62N�c#�bQO��U�}l��O��i��
Z��F�?/X	���}^��N����Fp�'S�_�1�n����V26���k5h㍐4T��ah��A�j9d2���R��� �~7V��W�/�\�X��S!o�؟�bՖ�rko�1�A���r$$��0HL#^%��R��!Z7���"bV�!�;a~�p�i/g[�:��ST [�hs��.}��q³��vor�d��J��P�L���`�K|��i	�Ж6!�m>��Y�,Y&�u���T���V2�����I�Ѧ��4T�e��E{�|ː�C�6�7������FV7aԠ��h�k��M�����%d��G�(��F����4��pw��%b�C"���$���viS�9t��|����0���A�I�&�"M�1U����s��Vњ+��꣸�2F=���:3��WC��ї$��"�"=�$�-��ļ,�qB5�B�v��Ms�I"��^�Ӭ���(Y��`�o�'�] vS�f#:���U��׿����z�l�(Xm�]���\����{D�ڃ�[d��v�r_P�e�_o��Ɨ7�{�������4�׌�3x�E>~|��7����"Ď�x�a�8��)}��4*�N��2���4��6��	�RO��������0+s	�?y��Y&�Т?��6+����:��]�-n>%J�`ܾ;�q>��#��K;�����^ڑ�#
r���zs�m�d�8�C�܏v3f�<���~<�H��!BXR�·��:bx!ۼd��.�қ����Ҡ��U�z���,m�깤 �w� �ewj�h�7���Џ�����-�v�K]�i�'8NN��^� q߃��.DK�:}� 1��S�E��ط��k��3������O��%���jZ�c�K�͝"����H��!���Z8�R��4R�W�
gR�?Sx�ts������ؘ�W��'v%Wq $#W�(ϊi�z�$�m�w.�"��۸��l hq�h���,Im������M���A�t�jj�4H��r�|��$t��&�W{Q���XGa��m)A}��\S����m|r� �����H�q�B���/�T���p�$qm�J��u�1C����aw#�e˻�x�-ͯ�N��c�_r�Tk����լ-J���#j�_�ul\$&�����>����\p	7���;�+=�ESg�����XΓ�>��ެ{��N7��V1[J���	A�cXS� �ۋw�ώ�j� �\R�^L� �ׂ����M�D�|v�猤�(��t��5iNl,����@tUYP)�'�o���	ZQ����䶩�k���4�Y�殰"�����p�b��4<�pV/՛}�s���QE=�d��v��=�"�3B��iy���;��I�rA4&�
��N