XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��͏�B����x�0���QZ�}\�:l�Ň���X>�xXX��}�=��Fe1���H�u^|�PB\��h�k�DNؑ+�.m��BMLܐ�����XW��N�B�+�Jg]��X�j,\}7("<�Eo�3A�'� �P{���|C"�^������=����K؄��{�<��o���+�U3�<�!=r���`vҚ@�Ũux�Yv�ɳ�AK>���,"�N�W�Z,�`޽�Hzmlڑ@��A��o�MÕMvV�U9����S�2ʲ;,H*�k�dn?���T�{�咯~!I�%���a�P��� $[s�V�n���hr���8�O���9���"%I�w�|o����쵫@�:N�9_]p<P�jf�)���mn��w�t��f���VQE8��:������E9S&]�����q&��Q����y7���[�+�u��3 4����6�/SF��8��k���=�0��b0[3r9*J�Q	bY�-^��DSJ�7B�y%E��vr����$d&W�\%�F �Q
�U�z�a>$EoSV�׀���X�܌��߳I��/��g�hM=>?PO�P����83C�GxM	
�\!~�Vo���X7��j�Sg��(��L��:� �J�c9/-~���(_'U�D�3��a2G���Z#��o	CtR�Z��U�,F�K@MW��Ξ���!7���L��ZR�hĳ��<c�D9���6ׯ@1 ���O.�S�a��ې(���.�!"��府�9R&�����M�vXlxVHYEB    285e     970?H�W1��s�g2�	 ��I����b��V���g�î6]���}j�Ш�(�5J�&Cڀ �������!��j����n��8�U8�y��y�t��Et:�{@��)��b�fj�O�&����N�]���)M�X���/�:�H*Ե=����|Û�ʗEV�S}�x��ۆ��jq�R2>�n�.d�S����P^���ǁK6)!���J�8;͡zaA��1�e�� S�"M]p��F�f�/�=⮳wk�y0�^����f	I��soP;j�K@�Ƚ�y�[>O�*�:�I]�̬���d\���?�%�b����hJ�4�n1��0�p�a<ϳ~	yd=���Yn;����g۝]^�?���FE�Uy���R]1��OvN�	�f�YJ�G�6 ';�1}v��S���cx£|*��t��!W2���^���Ziw�����ˍ�� �Q�76fQ�����
���#HN)1-n'�"xVo`t�|�8Z���¤C�ڤ��x0�A�2%���%q���u�I�o�l�~�na�Y�E��@�BQ�-o�[Nޜ!��?�pE"�/�2\�q��C�^�����-�-��G�� @ca�`&AKT����	��n�c�mZ����u`��3J��4�#@Qp�2�`Շեs���Yk��Q�es:$>�{�Nz��I�G�g#vs / z��^�1���'���k�4vVX���+����'Ϛ.��E�i��8��E;���*�Ì��,�p���0�QJ�ҍBR�?�\�F`�t�<Z��Z��0��z��y#��@��~?}���T�ڲ���{S�������/���pst�'d���$�*E�����d
V�4eq�袈1�R|��aiY8i�ڌ�S(��6�J@xF{���8��Z_Y�σ>d��e�;�Tf���eޔ�'��펵̕.��c�g}Z�W�>��[����?��؝�GM��G�	*_N�����/Z��D�4V�����,䶂��pR�칣<�a!9�����Sz�Pp��3G��y�����g��(��Sflv��IAw1q�'GI����R����*C~��pR�;}�������mט�Y�.-R��Ԁ}�DŤ��|M�G5 �}��`��~�e������Rd͝���Z� 0c�����JϷP �L˒�3-瑬���f.F\��)�N5
�<��S�;��:KQt��n�*�ب��71� 1�����7��R��D����񜉈_�qQ7fC7F�	���x��D=��}"(��2�
����fa%1�t�t ?�ێqŽ:�&���{�0w�]�t�h ;@�r���mK�{�9�݇Q����(ES�MW�1S����dZg��N��F�>(�2��YXl_PhN�P^x�^GA��74���G2����:��1��.V�y��퉇��69}��/l!�~ʚ}9em�|B���Y��8�Ƞ���k�-A{����\�U� D�+B5�����0,�ߡ�#mw�AU�:�~��� q��D<�a��C/��X{�]�xV�t5�fF7����5�SJL ��ZDl��9�,��R�	��9.�߃��sx<����R��j�9�/�;j74�ʻ��a5�{㼊q�~�EQ�������i
�5$�>n�(M�}8�Gzt� �ص.,���o�+V�UY��!P�2����OI��V��	}4"y��>w�&�o��l�86Gn㨗��-�#�'2Dm̥��XB^ӌ�[�a�M��q��;"�ݳZa2��v$�2����M~Br��9�1ݟ�A���;4�&B��g,y(K���oΌe���L�}�y��J|z퓂	�S4~�C��2g�|��6U��5h��o2sp��I��8u�r�kQ��E�����/�󍘨_��7Ȱr��7��6����������l���
��FL�1�1�̺��#g�ؼ��;7������u�c<x�龭����71�@�4����a�h�h~����SܓM�AAɖ0�%H����8�RZr<��]}�6�3�� ��/�R�\Y��jɾ�]V�H��<�q� ��D�9A�����X=gW��%w{� ��eI�ϲ��*zs�?.ȉ�>��[b0q�j�m�$ ���>�ע,�X�h�r`�q����i[ްj�� �pH�D@<@�-��)bP�.I���!/���G�CN�0�Mb��������֣̊��UY�|����;��|�Q���\%����;"�� �X����o+nZ醁�L�(����m^��aP��>"��v7O:�?俗}�"O �GJ��2�J��* ���q�-����<w"��\ ��[�f|n:~��}1��1c�ȕ�]<}�� ���Z�!(�ۆз�d�6�rt:i�0W�V��awV[�$