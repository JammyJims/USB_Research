XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D9��dt�F V3{��DQ�ﹼv߼/b)��0�0��r��ϰ�6��#��z
%�fg˒�Bo���fzH!�0\G��\��/0лj�`G���S*�^�E�����F�%wA*�:Z?N����D1y�� �Ѓ�!DX�D��=�xe�ҁu֧���~f;�T�W%�%�h��ͷ�*��*nA�E&5la��K)OIF�~������|�K�aΣ�)�� �ڡ�����^#4�Jr)��V�{���w���Q�^�+C�5�/ki�6t����ز	Y��dϺCT<���8iH&u�i�m�L@��\ �x����Dȼ���i��x���k^Z�yL^N���k(i;��i};��<%�k7 l�Aˎ���*w֎�[��E����U���x��DG��/5lp�)���V�rV���P�	C�b �Vw<舋o�S[,�yE�Ż�[�2j;�7Ѵ�����x���R�]�	�N���>-#|?=����/���'<9�%�ac��y�`�T��?�� .F�f$��� Q�
�����~��َQ]�αg#~Q'�r"S�S�+b[������Rf;Z,G� 6^��WE`�ۺ�=����q��8i�}[��r���T_$��D���hH��/��S�����>a�h��	Q���Y�-_A��w��������i�2�qv��8QF��k������F��Зt�T�dF'T|C""�w#�M2Ie�8�r�^��X�.�_A�\�c�?^CÖ�DXLo߼؁�gT�|U���XlxVHYEB    8c6b    1e50�}�k:���ɵ��Qv	�G�.˱�������E�QsJ��-趢�)��W�/6�Kr�>�v�+7���Z�#b�-�}�B\�7��~�7�I-TORY���0���Z��p�����@F�:>�-���WG�xĻ��|������E֬�mI�=4n�#MG$/:%S��4��e&\�j����#R���k�h�w���&��톫�^q��/N�`"�uˁV��)-�=ך��9=zY1W��8TG���|铩�ɝg�O�\{<=�RH�r���FC3��� .�p tèz�]�Ds�T8�ڠ�?y`>��;���=O��D,�u�`�z+��ɬI;�����f�9Qvh�C����2�u�2R� �ֳ��\�����AN�h1�Dū�H(��(�J�̒����!�YE2G8�u���Ae�Õ7���0�q�_.Ժ%ţ;<������#��ӪtSJZV�U�NN�/=�ｪX��Wu�0p��]��c��3!�-�Y�H���HӃʛ�ߢꡦ�a�5=bm�j� �0�E�ͱY��a�A#E��%���t`��їI����^����7���l?�@Tl��2{�3�5�gx�5I|%�wY6)Y)S38����]�1���" ���꘬p+ y�Cd=L�]��'�7Lwγ���	�S��13�k���� �' ���N`�t�L"#�g�WT���\J�#�1m��a��Vp4�2�~ţm��~,�tD�����H�BnÁY�)��\1p���D�H2��^��M��H D���Wq�]!�13���*ڎ�e`�e%��qI�j6?�1��ZO-�Ă���� 'J��5�b`�L��`�u������r
��ƹŀW�2�R��w�˝`Dt����|��f��I,1��*-/�p�!�=�� �}}���eP��bgWE�� ��>���l��b#���
I��pr7YU �gx�jYF!��N�i�uW��c>=��d\�fP���1��ʠ�ZN'Y���P��G��|=|�(3�PUք��F���N�wJA�{m�ƀ��-����Lfk��+ҹSߔ��`���{��5�F�|ܒ��[r-T�8�2Y�<�s���hM���Ԙ���bg4����h�o@�13~��,Ho���d�A3Iހ����!5�6�B��>x�0��<�`���g	~1z��xN����S����뚜�0=�IF��{�uǥn�x�
A@����knҕ�9;U`j<��y�F����>VȜP:T ��=g8�����Ҫ�<�����ų :�+-8�:��8�'���Y�Ix�K�%�/>���ekuWc^�ȡ��	�D=�h׀�+� ���:F}�$7(Z��%�St��F�
`��$+�F9�Y�]V�.A�3t�C���N�t���I��k�R鱳�
3�ȱ-$ �H�>�p�Ǧ囃f�fE^�x<I�c��k;&�H��t߀o�d�"���/��\��.�کkn�	�ކE�)�_���m��!uy ������q�����~�y�ih����!ך�X���3�u`�>� v.pTMKe|4�.�x�]��YC��\r�T8P����{�5���[���w�ޑ!�N8�<��u~"�a��5H����CN!Kv����,pƺ��A���R�	i�zR��������TqrXEʣ����M@�?%�������3-���'�ڞ� 0���e�t�٪@�S����s�y�����*Dŝ�ڍ�[�I�h"��yK-���E�Ǎ��v7��s�^�:F�.��y�O��<�;��v7�G���A�� 	�-˷ޒ�6a�؜	�@	���`�n�ʨ(ݲד�fD=O9��]�'�:�gwxvPZ;~�F�Cd���M;��'��<>�W��O=�[���Kt�F+�צ��(���7a��]�/sT� ��'V�0�4��23Gu����t�>�_+= �i� �H#FStm�����WM �(�Ko�M�)�{Y+�n��:����� TQol~��ll̎���H�zi�����.?�A��j�@e��w_ey��Y���(>�7�>	�eؙ����t�G�'�+a��������@)5	ܭa� �ē?V�Fp��y��YQүFτ{��``�%�0��AK/+.���S�!�F��<; �[�L,�.A�$�����ȇ�"���x���j��l���{�{ψY�l~���?�4�x���z`���(�̓y��c��6{&E�@JMj�V�����Qx
/ vBcr����:a��')�4r���֊W����'���*_>/a�Z�I[���7�5�� �l7�񪰊����i��U991�e�$ӣ���3z���.^�&��Y�j��u!Xg !�Ŏ�B�q�S�+^�ב�h���5��}EQF���Pu��h�R`��3��!��%	i�P1Bl�M�G�H�t��e�Uͨ�l�0�>��T���Ҳ�����qP%�B#��Q�$�
C'��'��vq��q�ܾ�
���B�Dnà@�k^Y�pC͒��[�G�5��$��YaK&^`��A�ُ �Y�|\���:q��ˊ.|�C3u�#����	"�Bję[�Zt������N����{]��ai^A\J�X���D�p���N��-O&�'v� ԧ�kFވ�ǹ�*����@@��h�8��i��c����U_�n[(�C�s�6�6��\�_���Ċu��+��-�w����J@n;_;�}�qJH�$)Kt0�w�sȻ��YZ���s���"�u�Y�b�~"n;�.@�}@�5�m[��jpol�#�'��ؗE��������ǉ���E$�|��v�x}s9�]-�ԟ��y�~�9S�2�c��)�P�
��M������U� ���s��~X��*䴃p����`eJ�^a7ě=�J���:�e��/��إ�sە��osc��1�	@ȁ.1�����zD�	ظ*-� ���;�j*T=�����l49'E�=���_L2υ�G`]�]�|��&�`3C���H�ƆN�@�Y�U���H�J�[Y�tr*�&�C*�
z�`�����+��o������L��7uŬ�� ���x	��P888<̶N	7t�Z��!г��c��,��27�?�rL�����4��O��{���E��l��g������2�k�O4ށ|�_�z�Kr�»�}�����i�)��	��oV̱1�b��9A(�a(��D>�&�qQ �{XR��^��-��>�6��d��lʋVu3!��Yc����W��۠�"�VQ��_� M�J�Z�rV.7���.���� X8�B���`d��k]m40e6Y��P+����İ��{⹹/�r��M95�m������oyf'��'ǂW��b)�<l��e<�o��i�	''Q9Η���o�9j�U�����x^��V�,���s��;�X��uA9�nnpL�>rf�њ���ɝ��|�I5���H� &(�s��R؄��w���JY\q�?q=a�y��z],��/������;J-�g������m\��iV�۲�`J�St�� ^�4�	�Q~�)jf>o�:/�O:'O��k� �G
\��0i��
?��?��-�njK�S�Y�����]V�k:he��,���tG{��j�-�����}]x�������T t��-mo�9?ܦ�mi/;��g&�Aa�e]r�9�©p/+* �:�)�Vh!r8�� j��^>����X�X|�j�ۜ]�Qˏ�q	�	����rm��;�ε�kȜz���{�Dz<�����g�^�4���O��	��H-�#z#�>�C�s�I��1� �q��ă(�O��7&��e���u�T�V�x�HY�<+5r���k�||ZF:�̓�0�|�\"�R�ڃ�:W<:��?�.��cC�#I/$�֗��)+�s"����!yrjO  �c�5�G8��}F�;Fg��d.Z�dN�;2#�d|�_���[xjC�]��~�l��:QX���i�"�~MN3��!�0�ݞ+P�`C0[W̜����;+6r�B}j�R;6���I��w��u8i�cF��z�=�.K��k��`C��w��BW�H=�y!��p��@}��p+Z�_v������X��vj^"b��3%.$0j�!����t��+A����G�),�J�c��(pM�yx2�6=��S�� �ܤa�FJ��v�ʘz.%�k��G_�wX�]����czx.)i7��?�3bb�$��D��7�*+�E��VX�
��b�r�`�����%�_�$�k��~��su<z��G-�qċ��@���U;jtm�}V�#����0�3C�bM .a�<��/_�;іx���έh�К�,���m�XT�����wAE?\�"�>?>��af6��ь]V�i%Efj�l��ݹc�l�G���7.����N�ݺz�b|apj=���2E��/䏢���ti��I6"�������c�!T��l���G<-�}����F��&&��g���5�Y�gϱ#��\_�%F�#�j]p�<�X��9#H>N�)P2ȁ*а�V�
t�Ru�	���Ţ}d�$�k�x�v>�At����:m}��胕YC�L�9RU�ӾR�{N߀����@�f�P S�*G�*_j7�+ ]�ƙ=�/�9��{q�Ѽ�1ο�H-�YC��ĺ�x��ח�=������/�>9A��${\>c���D==�N4��;�g�s}?m�9|���3>�^0�^���� ��NE��t�t�j�ˮA}V"���A6� �G�U��@ 5�!4��c B��G_���c���@�]�����г�h�q�Ê��)�����0���%�Y��o�����oٷ�`�E-*�w�{n��:���(��}����ch*�r,��9kj8K"�^�{"�'�+���V	�8��ߞJ�V�9H��fJ\���]+]�j�!ҚLw�|QY�Ƨ����Qx�����R��Fe�B5i[c}N�g@X9�r�CliE�JE�O�%8sN���\���F���d	z0X���X��1��������0������LqW��͙s�3�!���Z[Nt�p��e�k�];V�Y՗}��v��c�C�pk]��^z��H;k>oJL(9 m����c˓9L�Z��'b(5�l����.�GS���dŮ��	�k��w�Jh�3b����Bx����`���2.��N�@PB���ݹ5��ks���={�� q*���l�Do�*�D���
y"�n)N23�a)���sM;����d�s6��x�������n�-���: Ki���I�[���m}�Fy�(W�8w�u5#����Ɲ�ޫ7�����k%�C�C٠cS2��F��~ q��C&���R��K�0֨�+a���M�W�C��)l���H��Fɦ��*�kk�l�]� ��5��q�yޠ����O��E��C���h�>! �hE��4�K�
��p��tҬF$^����Ԡ4��]Må\�g�U�bY7����]3�Mt)+�M��_]���2x�$i����^%���I���o��i�Gq�d�|z��\_/Vj��]��;���9`���e� �AǖzQ�˭��>��K)w(��q_�~G!*nɼ)@�(��bRD��3'k�nW�S�m<����c�欒����G콛-q�J�����臘�!�w��Y�u�B�CE��Ć{iGq�b'��/O�kY��֛!B��?�� ��2�O�"i���=�ܜY/O}$�l�̈́�� L�'���m��?vRq�������e�w����ˮ���!��iIj��5�E��N0����e�Aߺ�x��tG�Y]ɤ�r�������a��ՙ>�[��5��-������B0A�Р[���롻�%�q��ɐ�$%���J�L\�G��~�)���;餺 {h�&A�T]�a½�n��ۚ`�1�s#-ue�����,����c�Х@R:��=��TT��B��}]��*���8���^fKJ����1�a�����^"���#V��+!�V�9��,��$Ң��cb�vh��8�.��i���z��?!�ۚ�JI�y�N���N��0�9�����"(VG���-��@�a�0b�܈i�b`d�h-���X�������t$�I�P�C�gz��T����ɞ[�G���S��z�Z�?>J���4EF��J�L�u��T������2�fl��4&�6 �; /�<�p��+�����\��D�;�wYh��X���H���y���s<(F|��	~j���!��/�3x�2��?��d�kok��/�����`v��El����}٭�@�o+�O��0�ɍ���m(��΀�� ȿIyR��3��F��GWP/I�!�m��H�{�����≴U��nuw�/�Y����t�w�K��s-v��v��;u�5�M|��}�ǰ�a_�"?N ��k�/�Ň�V�{��h�LP'dy�,.�I�H���3E�Ǥ��K\ܿ,�z��㈋�:A��$�D^�u?�n� �S�7}�w�R�q1NJ>M��/ѡ���%�i��k��IFq�j|�V{�aM�pMà�A���ै�X��3���|��b��.��������;�Q���c#4�}n����l�]/J��V0X�|l�*(fj6����Ba�-����x?P�s+�=з�=t�b}3d�-��Tb:n����'�<�ŏ$ �i�M(	̌���M���.9I+�P���8G˨��1�S�賕x�% w��E2��t�$���Os-����!���ލ��Ps@$C�%�)��?Zڪ*c�)�U��C�}̱i�I,�K�4���+F��}�v��W��h�
x����R�g���-ǂ����ޗ�^JWAq��ln�~�r�C��g�▇0��0VF��M=v����K�m"VzX�C�"�ZW���=�K�������-ױT���D� ����_�|�]�۲�;i|m���nN�~����;ρ�@u~c�*��"����?�t�($OM��r
�!�SJy���
֑8&Y�?6�h.�O�՟b�č����MU��M���F��%������Vt�ξ�	�~N��>�����PDK�=R<�
���*�Fk ��ُ���kt��1#es����=6'ф���`L�]�~��ydL�.�� �f�h���&B�lm���ցzoel�3>/J<+�o����^&Ӝ,�*�AO?Wtu}�ق�m�s����򆋵"h�	�P�WK���-��6����T������B�2gІ�K�2� �޾��/���k!��o���H����Q�:q^8����a
�?�w��P�ʖ�N;��v��nU7ʁ������WN����\�IK]�F(~�}����+�3��b�������KA�S=�4�D��Nҝ���kD;0RGt�pN��XIL���!ݠ�r^X%d�c�'���{��:]�ў�ɠ�g�`�"���Q��_�M�r+�u0!�\��0�we��������_q�և���ܑ�pE�˹"\����N�RDJ$|VԖ�mp�B��-õnZ�.���e�y�u=�w�_(a6�a��9zl#9}�a����A���K��
S@�<�&�4�_��u����1�nH �!H���?�^�*6��8֣%V���w��ݺؕ`�&�a1�j�5ḡ�:�]*#�s>lUy