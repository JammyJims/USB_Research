XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D��sJax8Z2����'��R�6�l��*3=�ٿ�ɋ�т��U���Z]|���{hR�["G��YS����T�T0�c�g�I�^�0x�N�U77c㩭���:�U�kw�m�r�fZ{L��~Iµ�K<�|b�S4�$>u��qf�NB}�I�uC�[���1����$�X�i�3����[Em0?(����ðe6��gG�?YbP~����HST���Lʆ�)�$��6T���ťV�N�����~ዴ�S$Ǜ��������N�s�"Y��h\�LJԔ�A��'��b�k���Ms3kX�+�fNŪ=԰/]M�V��~�9=�Ey���>�S9�]�c���e��\��i�W������^ؒ&��Q�<�1��Σ�.�ڏ�3[!��R��+�+q]��5��c�gz�׺��qy�GVZV��V?�nQ����{/I�Opp�(�G�hϽ��n�U+$Tl�H?�)��%��#��h���Ҙƨ��X҇�U�;S�x�r$0���$��彼�sN>��n��x���)\집���1�:-� K���cQ'Ɏa���
.�ۈ��_cn��ާ�a������2�Z�5nu�^�7������$�f3�&\[�m�
�.�Q�/�IӠ���	��Q�II�E�?n_k1�|�4�ڼT/&���9�=�?.w1Ai����k=�*Ӂb-�ۓ��>�w�cdc@�Q�w�!�F��P"���N!��9�e�I�%����XE�:^��XlxVHYEB    fa00    25b0rȮb���I�b�;��]O
Y �>)�n�	?�>�jI���9�v��%�	����Æ��
9L*��شc��]�O�(pJ� ���K�G��b����m]J�1B5$��}�xCb�f�Tzh3#>�Ja79ឬ=m��f��(�7�*aS��=ۄ�.)
^#"���t/�'�f|H�9D�/��yz[�4&ŔR�=�:�4���� ��񝣶��@k� I<��'�xӉ`e�O�4)�R��T�s����6Q	�r��J ��j��\�R�lW�[&�5�O�������X��e��/�!уw:��*��*�?����{�"��Nk�|N�A�0Ks���d��_?v}Av��d�U_�����q�,�%O���1@���xZ�O�E��X���T�Rm{pP�6���'���T�E�BHI��}T<,��j��~{OC�!����8����w� �MRi��%�n��`��3J�)+�(Wq*�CԗS�kD�`����dm3�|9��:�s�\MO2i��j]K�s��13�8[	O-x|��-�#�ء� ���>�,��6����^���r��� �=�[P���T��YK޺�B��/GI1��4!��yy�P��8�D�&8��^����1!D�0�0��fG���A���Xnض�u��`�����������zau1深�]i��mxxi)�Ge�S%$h��30݈kR�^r*66U��'��i����M�+��qpԷ)���k���<�r{F�2X�;���	�)����9������dT[ U�зL'l�Ư��64-�X�O�^��赦�����;ƅ}�r �ƅ z���^
�����7*���e`}����'��:�ݸ
|W�6�	!)oД���a��FL6渤"_k�
�9��ߕF��E���WU^E����5�Z+�똘��e|<L�|oצ�KC#뤚��X�VSqw.�A�SO�
�#2)��-��~ {��@4�'+ �����:�~�j�;�[R�y�C(�_a	n��8	�ϧ%c¨GS��Jl;�BY&�}�}�IS�]D)"�,y+����+��I��B0c�ua��d��U�6}����=�;B����Ëy��n�"zHG��H��l
��8Ze>念���W+�H��[;"E�� �j�%��$05����!��L��h3eg�1T�`
���hqoz��L:j�ib���c3�������:�Ņ����%`Ė���@�Y���X2�,g
P>K�/uuV�6��'�zь�����F�T��WrBv .���.+��3�a+H�AS�V�� 9����"?��U(���]���Zt����ߥ\��Ga�M�+vM6#��3��n�عW����f$Rf���'E�+؛�C�p��<ߙ�������g�q�KG�X�C-,2��#�7�Y)�v��B��pK��D���I�qR���?�k�.`iI�BX�jl����8�\g�g�	���vЏ'�/���8MM[ư&Y_�n
���<�0$���ki��p#Zq˫����VN�I+߫P�m6<sC/3�fl�$�t7��ɐ6s�L*�����<Tɟ������<���,��" y�`K��!mx���M������ئԥ3��X���.�%c���Qy��@���3h�ouH����F$��!`;�G����P�xty5̾a�H�h>ݹ��f�V�ܭC�3X�'�UB�/������!]���Vo�G�ŝ���*��n������j�vLp�]-���/�os��P/���Hh[Í�&=;�?��O�'���ކ��ʘ�<��3Ϣ��mD�/��s)H�$a�'�4�r-���5��_�����.�vc!O��@��G�&s������[��Ɉ�b"�`!sy�ҿ(����\�����[DJ2�q��'����fu^N��ԃ5���%�{Q�J�O�p�wa������ʓ������a�D\]���Pq��v�8➄�R+��/T�kU�X�K��W�c�&	]�7ۨ�1�m�����u2R柳s#�����E�j/����xO���@�ʘ�n�$7p[5hiJ��5>�5�cV�j�K�T����p�&��%�p��)7u��t7LZH���'x�e����:ƺ���xeam�ȹ��2q�Ms N3��CX���mh��M] Xcj�Y�L�:���F�s7��>��� �ja@<_Y��Y�Q�R�f0)}j�z���ё�V��z�Axm��ԓ�#��}�������WU9���U�kW��n�y��l���P�KҘ����l�u��7��d�������%ο_-�^Z��M��d�%"�s*�o�p�@��ȥ	�}�Zr9VG/ƀc�6#s��Z���������g�e��$�-~(�j-γ�G����[��l�a+�*�R���(��+L�yQ؁0G�0��H��^�v�=63}5�9�l�+w 2��8��n6M�"6�1g�9ytM���-䪿�5��
ϼY���-9�0���z]G��֠��M�����L���:5pYpc]�|f�&k�u�@R����MPwp����_���0�U�D_��)��+����\��B�Ӕ�i�q3���F���^<�E�+��gB��d:�Nb�BAj�-B�ī���\��$2@��\��г�Q��_$��@v��N��d���-JL.T�6Ӽ� ��	?����i���F�͏>,w|i'k\x�t��b�c͋sV���h�����,-tL����W�yght$�v��6��#8��⷟���sJ����>Y�W�ĥ5�:m��44�t��'�;a��렬 �ԅb�֒�GY$ׇG�f&綧��#��	ͼl�:��R�[�D�n܎ܨ�'*��&i���9�V������� /4����e�Ɂ(D��o�����M����=��?�Og��]��3I ԲͮGa2U�����.�/dVA��̞�Y�i�B�_wp�e���$�1X���j&�~��K2��߫�8?�h��+f�5�a;�\�� ���X}�<�ٙn�E,�]�d�eXm�blTAb��gzo���ͳ��#����E�{7r}��R:,���t��fQ�bxe��²	_�>��t��s��(wZ�hs߭�_,�)x]�>j%]D�>|�����p�>�I}��8�� 89B��/�UϏ�ya}��t<_z�,�*z�`#��?9��k[�q^��V�?�9�=�;m/�o��."���	F�u�pU��lP·R�+�"����������l��P�Op9����������bT3�ǟ����=�$��e�#w�d�Eqx�R?��1�$��Ro�k�Y�%8�A?hig�d�Dw6���
^��7j@��:��i%d���[�ߦ/(�x��5�8��L��9b&���4<G!-��[|a��Q�(�p�-��<j3q�񶾵l�#c�?���@��j�r�!�?�A'�I(iF	�\7ڬ��	+���yQ��qZ�}���Čt�E�_�4��#�����@�8c�X_� �.�;_!*�+UϻW��i5%XuZ5�F�z�r"r����z�O{4�S�5������5̌Q<R�K�n��`�CY�!�	���P��5���|�W�����o+dZ�ʅ���L��u�?��R��eY>*rNݼxO��Q��H7T�9��[A.�3�R�/x�Y���1�qj�E�JH�Չ�7�^�Ȁ��P�%��������-�fCh�Eٹ�<*�i�%�>i\B��T��l��x?�8��J 
~r�3G9�T��9pL;uNX�/�vu��-VTo��c�W8(�Vdn ��t ����ŊqV,��8ý\G��F�+���}���`��կ�U��^=��#'�z����́����l����GE����[}��K�����;�@a�0�GfcN�rm�F�X(�?�G⻸a�|_y3� 0zM��ˉ6����Rb/둗���/rk������x������š9ul�H�s�J���HA��)2�	��W.� �Q}��RS�2�G袭+���iֈ�zVN�.�B	̈́&�e��:�Hח���KX�V�?��O܃�jK��\��e��������ټ���$}��öf�
���Qܱk7�|5���W�y��k�(���m�H���T�������U#a�*L��س��w�.QJ����p�A����{<��\5��M�FؗC,�wy�n�-�`�51������*��X�t&����X|��y��&����z��xOG��4���r����.�
�v���� ��:�)3�����5%�W��w�:���uv�}.�ٱo䓳��[w�I���ԭ���0��O�Hƛ_Q�	����Qfi��b���T���EY�壢�~���={�.SA�#
�ˉ�7�t��с��q�4�_��̖_K`7��Y�E���F�������S^�C�ž��kQ=ar��\�+��Ї�jW|�W��?R�0���#����3�Q+�̄�]��v�B�Vô�95jB���O���,C��H1M��7�Q�ٵ��s6�^'�9����/��i��)�������iI;N������M�\Q�2(���.���`�p�5O5;�A��S��c��Nz�#�����ŔYX�Q���>6Gq��}Wؤ(z�n�a[-i��^(F����1cY����3���)�O��$]�qu�ɚ�X���Y�_�f�S.���_�q�خإ��y��y1{��\C�b���ql.tF�Ӓ��W�5�"��)C+���<8�����r����1���d�x�W�a1��,� �u@ŵ�2�_�h6�W��qV�94�i��\�d�G{���0�F���K(SXaIۺ�0��:��d���Ox�y��s�;H�#4\Ʈ�}�͉9�"�*\`p��Ǒt��%
2B�X������Ν�L�.KLP��:8ݠ� �.�F����5A��8�����3ɐ���~��< ;<1X��xJ��Ѫ��w��+n3A�|?s���.�w_|�H;�a0� &YPz�%K+p��g&6��y���`3IT��p��E��&	/we=I����`w�Ǚ�<�S��]$0M�8� s���4o�	��Rv�jD��f��D�ɶ6�,m�x����uNGȑ���f ��@ 28�6v֣>8/��Q��h��X�=I�6�%2z�.�zӺd������1+��Ӳ��;�fM�f4H�g� �`Vn�+;Ϧj���
g��N;9g�d
�0�R���<���J���0%2�&�v!^�M��C�QId�cwױ]�+����h��U�[�_n�S��=���+�%�{�S,(�4�2���߷%�aMؿC���܏��
w��oqh�$(��O+K��X��|[?Y��f/��ǽ���x�KH���ӏ�7@_���J.�{�E����^@=����A����0�?+s�� �6$��q�T�0�5����l�S�	��&F��EscB�7B@X:�>��
d��q~఼���A�s'.�)����([�Di����W�Fw�+0���V�2�o���ݚ�1O�G�%	�_�����+r�5Ej����
�� �A�&���+�qΩ�,@S�Q�sd�0�KHr2�P��w���@�ӝ�����R!GJ��B\f�<���V�W�sE�/_�j�	��WҦ��O�����x�ԏ����ʤ(�uIj��`��끓�d%����
�4|�i�bn���w �zK�s�о�s%dQ�oQ���א@~����*��݉Si'�p�F	��hf!��#����/���6t�.j�H~)#�����:������_��g>�9,e>�q�?��¾^���m	�61��B,���
R���8�]�Â�x��	�9�o�����Uqs��o9��FX��^i�O8m*��p�M��}m�?Mib�uh�@������R�ɾ�g�͡ERy5��@�\}�B��Ml��$m�d���qIoa㺇i�sz�Y&ҭ��1�&Ǆ��h+D��C	+^k@0��?���a|r��n��hr>e|�p��k�|��UHU�N|��my�x�YGD��*�V̌5%V��2 ���8x�p���\?9�����}��#�� �JAC�p�ч��vͯ-Ř�+,��e�FM�'��I�x-���0S��O��c�R��F��wHs5Q�#E#;������J͌�`�ǌàN�";�N���>���_��&�cs>���G��"Z��Gp@㙦nK��;K�#S$�۪`ΰ؋����'Q�Br6����Y]�u_
�BJo�L�fX?��w������֣7���U�'ҁ��ȧ�<��V�eEM����[I@����~���eb2���wD��N�W5�~~e�%^��.˿8#��5Qx��C�Q):�,u���7<2a+'�-Y�%3�XuHVvdb4b�8j��>��5�`I(�d)!����G���ue2\�Z ���ѹ��8�Z�P3r��PF�^6H�l٫Q�wRHB�FE)�d���&S*�@�2��5`/!�����C�����=ϖ�������ƕ!1�5x��/������L(�Pz��_� _�\8^S�[9����!f�`�Ɯ�F�40A��}`6��ר��an7:S��
����9Tن���#e��7%�)a����a�{x��V�x��E��ۡ?�뎺zT�,�=ڮ�9�V��t��zE��N��}�ҏ��rL[��m��Zl�����
H��(��e݁�.迦Ds�mz��D�U����8m_���������@X�lQ��4�5p"�1����>
���Yy.����zV�Z��|X�H�3v+���{��B!S1p�E/��8�0$����:=�"�_�s��a�HfbS؋%2�B؝�����uNI��_�9����Pmi�HO�,j���K*�I�}���?���;�J���?���l�YnA����Ȕ
�M���\��5���B���@Ϩ��'O46���'�[�-1Hz�27�P����C%�� +-h�{�>FuV&�e)�ᶔ�_r< Է������I��z#�Q��v�BK٤�E<'XZ�|�Ǣ*`�~
�o�Y���]"�R�Ȕq�����56F���0X5厽C�N9*��X��[�8$��ka�V�դ���x����8��Ɂ}�p攣���U������`f7�U�Q�ֈ�wD����)��$�����/S�ɰ�K�M��w0�;����|/B���K��v���"Auۤ��x�J8ǎ��X���L��
	��\g����8�g�W�����}��N�0Ў�x�{ݦ���2l�i�D��@�y�9B�RY�;$k��{5�%5���5��8�W}_uG��(���q�~�1��04N޿�%yZ�˃�.��)�\k2fYfHv)���_ژ2�:�����A��+(�b� 0z��L��J5dr?Sc�� qE��|�2�;{
!T��w�2&d�W?�j�v���L�ޯ�E��$ˮ��A����Q䟰)9��x���S���!ז��a?N��X�u��Ƣ1��{��V��J.QX?����XL���5���k���}�j�!e���cT��Dd��*�NYwo����i��o���Y���J�-�쁡 "�����cf�����_Qt@B�����d��_�׎��d;	R�F�*}TՍ��TjHЂ����8B�j��ᕗ�� �nF�8}z��� �^1R� �L�t�J;6T!Ϩ���ύ�zQBR��Ԩ׍�_���dShzN������P��Z����x�v��v�v�І{��¡+?�Q�����*��m�ʨ�4b�$Xz°4����L�+N�_[4�7JЈ�u�Qţi�UK����Cc7/=����}$�C`��Z4��MN7�K@J3����m����	k;�F��c��nq���kS��Bl+������~؛յ�����I����-e��5�a��ŏ��F�@PWbL4.>�R��	����&ڻ'��H���$�@����-�&<�����|\��ٸ�L�g^H3a+a`Ç��Ȩ�����k�}�f�L�F�A��UvQ�>����>�7쏂5Dl�R�`I�W��{_	ی�6r�RFy���|�D�ۣ"�;����a������E=:�wET��k��j��uW�(�:߻�x�r5w���� Pg]�jS�B��Z {�o�;G�� !V�Fr�}��w[|�@�����pah��-��44ځ���K�qU�a`R�Yo���+8-�+5
��⹲U�cJ�DO��ɇ/Rt��*>���������iN�Nx�D�qz� %�!1II�C�6�ieN��|�K�#w;N���$����֓LRHDY�<�i�6�1p�t�tr�5a�=>�4u+a$r@�!�����|���x2.y������M��"�pPi 0�_!%�ބk�=��ʯ�9�}%�((V�/��l������5��T[逃�/�Re@qzt�P��v/4��C3�|T��֣[�m��w��z�PE ����OZۦV�I�5�b��g�r��隄On���WaA��A��B��l�)r����:�(JFp����/,�߸a�La���b� �|�.����ɨ�袎�H7"Ln^lB��̈́�&f�A,Pb��Pw("���:rT�a(��i;��N��T��ŽHg��9���O�DJ��̫�w��d8\�9ϐB�|[_���	���FIP-�I0X���;��>��>L�	D$��}1:p��q�_��,�Z��I��,V)*��R�q���o\�R�*��	�3�}��&�1��nX�x��o-a���j��ʔ~�����S>~�����2���s�U(&WD���G������p�����+0g�?���MX����1���W��Z���G�׀/u7�n�]3��eK�ຜ��}����(�	�2�ӟE�t	��c(�*���C�4��2� 	�N�֊M2�[h�������8Sa�����"�I\S����^j $����!ҧƕ}���C������0ΝB�7���*I��S��|�� 	��~ψ���^�K�fIuч��SIw]��RF߃]?�� ��������`�,/3�@�r#kR�s����_��agO�5?հ�pw��&�k�~�a�>��&dP��������z=,�C������1�`>������ �}��RN�R9���V8?�=���{���F�5:���T����K
�\��������Y�{#�|�[��ɞ��(C�Am�N�� �҈���-��e�r��)Ƨ,JOUt�h�vP�j�$�i�MFu�NXCs¼�z��ǻ�@q����8�@�se
k�J��j�ඛq�H����c/$�$D���݋���J��0��ٗ?�@��+�x�r��z���e��OF]ز�0��n�����-J�mS0	�v�w���)t�p"W-�}W��7��b|,�E�i�i��!������J&��	r�{8XlxVHYEB    1de9     850XX�hg9��-uX�{�9cV	\�%n�(c+Û\�x0*l2nmww5,�O�k�D0�����SzW��EU& (G���t �ioZL+H��c;���U�K$��.��������0 �Q�F�|fa�'�`h>�����Su�1Y�w��M�1�դ����;��Ð���I2�V7�f��"72L�kGW9dꈕ���;�HTG'ʽ���3T�f��`J�f0�jqAs��;L�(���m�I�`�<uz��s��nu�i����2� �_�ߌ�7/$������.�FY�7��j�����^ƗH����J  T��nit.	�@�S�n�w��=� ��k_��n���>h�5���bѠQFwaO����`�w��l5��"a��;\��TBa�:�d9J=�����#��"�,��I�>���?
<��h�}����d�{}MYiD@�$	Y���}�5�����Mp�C`���6��G\�#�<���N�M�Əy�6�oq�E���/Ѱ�b ���5&S�
���c�f��0>���MM�Ȱ��_IB�ܭmWA�ߖق�͠ni�P袂�A�����*��R�l�2$G`.��h`���E���I.8#{ :��>!!�~���9ήl �ɵfT7�l��('��!��',1�v�q3}HB���j��b-U���H����ewS�2� �F�0fq_L1U��|� d)z���^�am[{h�zn��fb�J��RQ�W;٨Ħ��ev��P�*sv�����c\�.3"ma^�]�sm��Ge�B���o{�j���������z�����{�cfd���
	CX. &痺��Z�^0==@¦}g��b����*-w�����dg�5yn��ݜ�[�N�����ni�K:�Rq�d��]��5���D������˴���-=�Yf�g�$�=�	�@�z ��ǔ<��9L�1H�6��2G{�ĳ�.FoҶ,%<��e?*œ�]��q4(8�;�X䱔���DX�6������C?��Ę�G��P r\�6�7x�Bv�z�׭���V���7$�M�?Q�Z��`3���T!�w�����5a[o9;b�k����?��#A�Mt�讗_:^_�������i�a���(��2���v\��(�$ m����z�Ra+����tw�*���6E/��[���o�\<'�QG0'�LG*�n���O	�b_�2q���a3J���IA�k�Wɇ�f�1�3��t�:_��u�*�1C_a��r�)�W� J���3�H��S�=����ͻ�'��ya�q_=�a��M�&wQ�)c{��]�V�m���Fx.�Tg[������i
fP}�ve�d�,F�)��
/��"�1��V�A�Z�����gp�Y��{"�(l�瓩�mجn'�$J|K�B�}�,u���Ad[�6��3S*9q������C3�v�"��+_k��8=�7�]N����|e��/�������g�������z*�j���b����O�Ȧ��=�-Sd��}�i|@����o���V�Т��%�B�0)<�o�%6��dك4_eD��kzьmsYP�r�Bˠ{w�.Cl�Ĵ�,ף�\q�4[�u6u��4ͣ>h
���l��Z<��2�_�śbc�����:C&ψ�	�<�@���-hy�������^Cd� �G҃�_�!q�����r�INƞR�mBd������ϰ���!&{Њ�P5��k�	e!�Z�m��z"e*"JO�܌����o���{�rò6,=W=<�v�l9�HU���^���8�a�ظ�{�>� ڮ��`+��Ĕ��#�l�g��A?P^�\�3I�Y�:͗��l3����D��A�����>X���FJ��qڴ$�'���:���fW9���0P$#5��E�*/�ʳ�-���Zv~Ç.:L#V���/e�i%:rp�H$���OG��z��Ņ��r;8�`�]�F���Rǋ<�T"�jd��4p��5�b�����')�Gө��1��d}��#�l�d���
��t�i�k=�?ZEK�����s
g�a�}b���b����2�}�1^����\}O���-#��p`�ƱA��_|_��w�o��