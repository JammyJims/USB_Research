XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���-�Wd�}Fl��MkŅ�+���, I�wSrm��U0�w�]�5~V�k흑���j��mӮ#���gC#�.�����\���^��[�)T&g���p����r
�K��|B�@���>�]o=��|+vSE`B�����.e^륾=��O�J��ʇyj��%b
��I,Zt��	�XBY���Ʒ�����?�w�7ï���1�&9 ��=r�A�B�����\(����J'6��KEδ�o|�?@I��K���LJ����?��YA3���`���؁]1<%I��Z�旱8���"fq�K�p5������@_�ۦ��]�5&�;��z�.&��m�d)�
قX�Ip�G���QQ�Y�{�6�<'�
k��ʻ�d@�Q]����k?q�E��>��C�MJ/U�n/G�}��Q�'V��lj�뇥A�8x�H{;�vU�V�K��]�K0��<��  �K��o�!��Q�p��3s�/[_�5T��"p�yb���r����ޥ�C˥|�ºW�gi��@P\��S���6�b��b\&� ����~�,��FY6'e�+[(�q��=B�R/���s11{-,d|8��
���0�����I�i�*W�~;�i��E+2^I#�<�ԣ��J&Qp��O8ԅT�8P����S�ubW��)��ʾ�j��G.!b2�+�a�nEh8�f�(?#�D۶�a;@��@Og���3� ���v�{��CÜi���%�
��{Gj��9��<m���T�� ��+��cXlxVHYEB    fa00    2c40L��QB9�7>�^��?a���]A_����M ��*W�&��T>�K�g�E�cg��R�G'�yMe3��"�UF������H��J�JB��C����csT��s2�Ј��F��]󩶦����a]�Q�ƖJ�_	���F�l��c�P�>3���i2�9�Q
�b,	ߪ�,K6#�!��gε��)�C�����)�	�`<�E��"�]N&��V�#�E�
�$�FlǼbk��}H^��1~}�[N���A���\�����,�@���bx�uB��S�R�U�7������'�݅=|/a�e?�§�>�O��W���H٫��������aC��F$�7�b�V����ռ�Y��k���U\9�6�jc����a�wcQ�1�j|f�r�w�H�g�����A(~f/�O��滟KBn��pP\�Fpx�Fµ�Vg?aX3 ���p�#kb� Z2�x�������D��l*�&ՃXI� �~��Sh��X:�Y:3�ޭ�V<v��]�3=�	W�ʏw��3S5�*.ɭw��	�^����o����`����~��O��5��J��ѻ��T*8�$���8�Z���������,�?��o2MP���NSi�U %��O�������:����r|�7ne����+�(�gqM������|���b�R����\���E��_�qL�������Z�N��Dpԟyf����)֟�����l���ۤm������"s�4���}�//y�����ܵ��K�l������U�S�,i�=
����g�����+g)dLg��E.��6U^XS:���H +(B��ɫlcP�h�zII A���@n�� ���&��.����bf�t��^ӗ���o��x��Ye�����o���:���@_B�.N���$�؉� Eq��%��4�IdMf���+�Q�ؽ�kZ��M�h3k]��m/Fғ��v�=��W��Ix(��/���+�)P<���GW�-U<_����X
5��wEZR ��Ir�*)�& �:r;���=/%u�v��A�.\���4��t�{=3��3���j��^��6I��x�,��|��Aqk��Ԗ7�=c�Qz~q&� �?�k��!6'�8Z�%����R�DG�Pt�xO��#�A�d.GGR��!i;�?�|��$ V�A�?��<A@���̛֒D�G�fr��*FȔIdq�����e��h{���z
�A@��hz>jA]2�-fxͣn��o[���f=�Y�q)�@ãH[,�����Kǫ��L��&�_c�Wx��[����R�a*�g�@��*e�^� 4�zc�����U�0�D�_�:3�:O=5�	��+�M���1�Cj���5����u$j>:'ڎ/�\ƛ�b��<
�d���d7!������G�Ayܠ�J�,���$�(	�`�va�#^�-��X}���_��8���l0�����������h[�Ŝ��cðsS����J�EVl�m�[����Ob�ziC�M��x��	j�+O�(�T_ܲ&:��+��8r#"��M���s9����UI8Tj� ��K5��e��j��8�X0Fh8��P�W����(��ԇ��I�S�u4������mU@�,�X����D���ђ�w��Ű?ȇ�Ȼ �7R��>��@��n����=�)!O�hK��t!�������K�+���X	�:6�3V~������3T���eT�:���w��c����J{��~3 ��0��Ɉ��ȃ���
�t�\k����(Dw�*|�k:)��;��r�K�y�4�P`�Q�y �eH�H4u��5��ٔ郟��yS��>-d����)����:�>�ʢ.��l����h�w��h8$�����xBN�;X�^(��{����M��Vjw�t�i-E4T�m��Yw��=��//��l�ǿL�5B��YS96�������Jgr�`\^#tgg/�d���T��{]å��A�v��F4������疘�68��c�H�q���>	m�������o~v`�C�*#P�,��a���y·[S� �ߕ��(s]nCM�e<o%D�2�
�!\ �0 J�{�����c�bb��>�dHZ�����S�5�e=�uUS��K��L���@P�ڈ�Q�����OKQJ�~i�̑ߔ��D�f��J֙<VW-`�M@���.H^]��Zd���<���2�SK%��>;�,�w�9��Y��u_��d]�ז���l�ck�18HF��f>�����&T�	����`���yY����(�>"�^�ݸo�b����� ~��V�=~C��y�O	Č<J���|3�Q�x�Ȕ?>��72���c��8�{���T�}�27ΰ{YW�B��p*g�2����jZ���̊����?|4�(�'�� 	�w���{]��N ��m)aܹ [4P�"�y/�]`�L��
 �	��I~��[�T�=�RHƹjB���&=A��OT���%7�;!�Y�O�E��Sh�
�O���L��Q���@���Gg��9ʹH"�C�
Ӎ����&�j��a��M��-�N�r.|�,�4/t�%��AT85~��b ��S$$�����"XB����T��7`W��7/��M�~�Q4ؒ�:�,��Vvڸb[��sB�orKk�T�����s�Ze�z]�0�_�y8~��d}�1++|����K.7ki�:��-��N����%&e$�YoyL��U~v���:�X��S�����*jB}�P�p�"�'�d��W>d��z�)箭�T�����6\�6�>G��b�I,ƞ+ɚ^/�h�(EDM�Vdj#�����ZM�i�Eχ(g	�I	�(gi0q2<���}�R}7r��İ�dc�/�1<pq�;x���ì��B�B��J���t̃j#Q��8W]w&�Ø�g ��)	o�>�upc\]a�JҾ�CT�D��A�@y�۱��/S�*��ޅq
��klj�����r@����^���� )��P�L�O�: �վOA��AIkfǃ�`iH�a:�N>�^�V�<��q�'`i���
n�M0���{�N�%�>G� �$��A���=x~��@��_����T��܊]"���&�?�mV�^3[	򝈗n]�W�?--_�t�*v�Z�r���ޢr��q�xPII��Zޓy���z�n��nGP��Q�Lq�-K��M.����o�b���Wj�3�����d��^��:�����&�mm��h6��Q�@�y��-<X���ӑ��5�/ �Fc�q����m�ؒ;��ʩdJ�|P��������_�cBQQYH��hǅ=k}�ߍ	��]�^V��Mk���ڿ�.E"����W���Լk.Y_�#�E����x ���%gŚu�<Lu�,��I�A�PF��F52�iK�䀕O˥Z�!	�P��\-�Jѧ�����r��"�Ђs}�=� ƴ�ך�j�Ӷ�TM�!'k%��s��t��H�;\ijە���(�À�X)����;W�ir��%�D����*�������Iԏ�iYޅV����.�e�3�)!�X���8�ۂaצzt𙜐��7J�=yOv��-�+�F�ͱ��dQ��	%�\�9��ב+H�6�BK�QE�ed� m'#�~G�uyU|�4^/,�!����0���o����gϗVb����֌��;p��>*2��9+��ۀx5f6a��G�h�P���K��<"~ڤ���tXlkIM��ʂ���z��R�#��t,��
��z*��u������~����?y�ŮY�<�>"��y���$���`#[�#��?�}�Gq�r�GI6�1�it>�D� �3I ������n�y�lHj����b�%�)�;"+F���:{ˤ�X�x�����Y=���}�e/#,羰�V��R�_���S��~y[�8?/I~Y��=y%�Rқ��v9�w�y�s�%S���Lp�^ �z�a�opҒ=��jm���t�*]]���,n��6JF �6�p��`���2H�` L�}3�GT)���O����\�"�v/��ѹ�n証�{�a��	��Jh ���#�����֭%��1��갚�\"����� ��'_���w������܈М<V�e�W�!��l�)�������3Q���Ro����'<F$:��]�!��	�R�Xd6���ڣM�|D�4��H�I����71��%��]^�~4fi<qq���(9�aN���t����C�.�ʷ��0���t���I'L��y�Fs�R��^so6�O��`����*���Jȋ�.�L�a�.Cu�������P�=��Ǉ�%��W��C����@$TObrJ8U�,�pW�Z�T͆��>��a\y��Ag{�tN���8F��q�����ϳ�v�%U-����[rD�y��U^̗s��v�7���=���N��`��0��S#
i���.9kbTL!⇲���7=��C2�V���'G�q�v��^�3��v�W���k�c�_��nN$����"�]P�W��J�Ʃ�3��
�J�W��U����usz�ꩊ�N��g',~�@ M 5y��^U. �
]Q�����N��jw�:��4|��َZ�Kv��3w[��m�Xp�E���W9_�o���g|M�s�#����♶�ׂ5�8I���7��y�{���~�:���ZZ�� ci��`qo o^��o\u�s��l��N��w��Kv֧�Y(��^RB�@$�v����y��w_mxmrIٸ=ْ�ˈ�����F��'�[�܊y��z�ځ�'z��|��R�{����NZ�q��p1�
';^;�䬙�¡�=��L7��9�op�ݷ&EtGƆ*P���Ͼ�YX��_��j��*�!��ZA���Ĥ0
�o�β�7����o��$�4�ld^��d���{(���H5OhB�����<��V}�����6�Ƚ����,4��?f/�����5>EF c�ו�s;�����Ǐt���yc�T`r���j���I$��6�!^�i�tb,_���%�1�5�N]&A}��T��2���f��Q$'�g+��M�jG}��op$n`UД30�}�PX�W�?���_=;�:e��+�:PW�ӿ��F�<�h>�U�Yp2�:�9h��mH���bB6���Z�"l�ڗ�^���R�.��(+�Q۴!�-�t�$t9,��ϭ������<O`��聉����~�4�2=��V@u{���K�6�N����׆fD��׵66�,}����N��h�l�fs6Ț�S	tn��$�����]�@�M�I�"���K����Q��Ȝ�
���?������Y���hħV�r�����Z�=������4��#%���j{M���i'�60��V�&f�3n��'�Z�p�ߴh��Ҥ4�ef:��Οi����ig\�� O���h�2���#Y��4nɫ�o7�]�v�y�EG+������q%�`Gq����
�7�)����H����'#����� �#���7}�ȿ{�*ҙ*ɾܷC�́�9礞���A>=�P�Ac4��V����� mA<B���^����h�U���� ��R�[�n�oָ~9���Ė��<���J.�$�{$~���������U��c���K���fqa�`��v�d#PF�L���q_�Y0����&��42"|Q�*��l�R
�L�>���U�`���U��.����RW�&6��w�`��=�
ل&��&ܢ����/)��[#7	�ٳ�J�*��ZMGK���|�*hTU�􁍈8��o�'�; ����%v3䊑�ŧ�VH�����V}'�?��&\��3!ʐ��e7f-�8��h�:C�Ӓ�+Qs�03����������r�=Y^)�K�&�6�E
v%� �+�1�n>�Qy\������o(=?��Sdؗy6�M3jC3� �:�����Z�ol��6�L$�sk��R��A���Oi6ɵ�L�P��~g7Z�lR�c����"�\͘`� n�:F�@�.T);���oHt�Su4ܖ���h3�q�/s��^w���_�L }�ƌ�3Z�^zv��a�kRW��2������L�4Q�b�4���a����D*�Q�uWlJ�Cx�X×�M��A7Xc̃�����M �C-׊�����]��!XX"����굕���V�3�.�z��5�H������f��KYw)Mo����IY	��PS���&$���}�o�M�sm�R�>a`�[�ıb�W
��r��`͛�A�-:���Q3����G��{���w"z��
��X<}�{�Шa�C9?�XZ@��?�pJ��Panp1Tue-�(���6}�."�L�u�pP`�q�����1�-��sk[�(���	�#`��3�N�ӻ^�7�%ߞ'x\�K��t�H�i�`���-�\�"=:[q���m�%��X��ܽ�p��e%���Dsc��"�Ï����Ye?��vm��}��U,S���K�2m�6_'"�h��,�T�폒 	�D�)�Q�tj ;YZJ�R%<��q�?�y�E�lZ��ȏ79�m�^���ɕ�j��רx�*i�C�<���"Ijt��oֆ���(���-yҐ���f�<���I&3$��P)G�퓭�M�ZD	�k��J��#PJ�C�5�I������i	� �?���B�O���=���˸p��%��+���qANQes�o�$^cp��.b���4نd�<�<���)ޠ��3��X�ʞ����H�n�<�p=�~�Bٲ�m1Ske���
�\�"�?�"����&[���|��K��-V`�g's�K��6rz��Y�\�pnȌ~A�
D60���cr<��hUw���(�Ѭ��Pl�l����q���ѷ����x�^� �zq؊A��������$��G��I�l=)2z���K͠J����Ⴧ[]����\�A�
'厘a6�=���}��U�5�'PcV�:�_�^w�ߑXź���9ּ�����+�7��~��=7X�`X�fR��L �H�C�dE�R�"_)�����f��'���%�n*�*E��8�Oޘ�x}���A����(G�q(\��(�Y�Ae�XA�X���(n��#�V�0�ł�h5�)�.c�U|E`�>���!�l�E4�m*�9��ʁq��D���A��
���|�ԓ��FU��9G�޾��We��T��-���y��&X�fU��������2^�v~���G6#��9�����>)�(=^�am\q�_~������JQڑ���2v��<]�2���ϴ@���A9�P
�	04,K�6})X��'��øE�⬟�"��(@�J�[5�H픹��ʲ'���A�����@!Dp�1�%���b��?���M�4=�ǾV.��k�?P�uK��遍h���l�3��
P���Yn;^���Lc]�Qle@B��!H=�rV�H@$%ң���ˤ#R���3��D���zpF��#���!&~>��0�&]��0k�4�(�)�S�p��i�Hԙյ�\��2#�/�>�b����q}s+��zH�Sw��Н��j��]>X��Ā5��~H���j�\=>��%��B�!� dʯ����9Ҟg.��K�lkL�U��p8�OvτD�L�~�����F�E1|v޳��
1��i���6���P�L|�����?��S��0x�C���%+�\�����V�� ��q�^&�*�H��Ѯ��6�?�ې ��I�3Ў�X��,�r>Mθ��Eζ�������)�6�d�L��fa[ޭyH�޻{���[���ʹ\>X�g��_h�9!^�Ey��l����0��z���"M�S2�5s#����@�pY������W�v�K(^�����=��r	�n��Uc�{<��f����<$����e�Q�B �Jp9?=�`vn�񒹷�IZ�]���/K�x�*������I�4x���M�#���r���9;W��F�<pì�x�l��
���j2˺o�ZkI�߲s�9��8^�B?��q��HD�zǕn�d���y֣F -�����Fn�%J���|Ǐ���M�Z�71�A���+�1w�_����8erJm#�q����Z_\�	��x�7���"Z� �g���ޟW)����~H��݈k/Ϩ���p��xv~>PN/��b�Fy�G��$*&��dv"�d5��gҤ�[��Q���ݏ��(SK|d��h�y���b�}�O�0��oA�ԽJؕ���}n)��X��^�-��Y�㓝��p�y7`i���n��&��2�~����3P������{YAc�R�4K�^����+��O�O7w��Df;�	����{]CQ�Bb]0c�C $��E����}+o����m	�U�
^�W<_&��!�-;�p\`�� |A�ۼ�y �{�0w:,�s_i>O_/֒��_Y07�a�B?�2��g�U`�ѳ(l˙@�>Vf�Q'+9*(<���K���.��1ynS�j���=�փ+KA?���ңޱ�;hͽ�>ph�t臦jɦ��<�1B�Lhf��P��=�����.��[� ���I�2�9�K/�-Sss�8ʚ��ۈ���Ҩe����e"T�n�1>b�����4����l�e�	qo��s���l{%�*O�A`da�n�?,��6=� S{��}lz�{o��C�I��PKjA����Puf������1��K�����s��7�ٖv�ms"��L�3M�Q��9�� �p�ͦ$+ML��ج��w�cc�8���ԡptIE]�_?qX��]�~�d=�����A=#�$4q�n��]��3F��Ѥ����1��rY&���"�9Dj]+�Q�c��'���5p8��T�n�`p��_|Bd*b�2%N��߃�(�wjA����G�����_~����E�@�c0�d~����y'*k��{�10�ڌ�KJ]�	7iF��]>\�v�/��4�����aY�!hF�Cr=�z}��8��;��.W�V�S���M��J3�v��"���$�V0U�A��[����u>�͢R�?�]i0e��e��x�7��TS2�n7����mA���JXF�{��z��ھ�y�[4n;|:�/FxW�B��P��#�ghz��H�BQ� Օ~�1�!j��91򓚄:�K���W�hEX4��\�L>����f�)Yd��""�
��[�^
�ܵ�H�U6�X��b���0�ߘ����� �>'�m���g�f�
 +�֘�%oi�EZ�O2��sG`IRް���hyJ�1Y�m#wm
�=3!eq�w|i�6��=���cQ��{Ϩ"U��Tȧ��Ͻ�� ��t�7E*�"O3�bi���A��/��u��٤�&{��5E* }�}��\�V%��'��2�����՗"S]5&�s���1�l�*��ȸ�C�K�>��K���$��ᾖ6�� �"�ngt�ȸ6���p�ՌJ63�!Q.���}���V��t��u���}���Vt��x(�V0LmxO��b"�;Wg��$Y�;(ju����1��̆���38�r8���-�ϛ�݌�����5%������`�H���q]U����Dg�B~/�����b4s���"S�`��F�C���,xh�Ѝ�袩O��e�-����+�$��`�1�A��6I�p4����!Z�.IKGE8?�rz��r���66�":X8�i�I�����eȇM�oӜ���6�C���Y���4�� B�zp:b�1��!>H�C.'�o�c����]���Y�?�$6B��U� z'FR|M;!"��^9��i������\ �O�߃�M� ��Od�̚�v����t��Z_�C�x��L����C��֊A�Z�c[�(RZ����K̰��g���vnt��=�F�η���!w�.�X�*,JQ��J��G�ZIg��-�t[�_�)f�0뵍[�H�.%�.���D(�����=2��n�+���d�zdV�2KJe{��rh\�}�X?9;�]R��"�sR�b�Ъ�h�rC�qo>s�eH�~��1�Zq�G5���e Y�B� � @
�[�I�ם�h�K>��h*�W�w����F4���9[ʮ�����t�B	dRw�%�3��r ���CBdE5���>���94��a��,����}��>=oN�Ć)�9�E�{n�<���$�ޘ2e�;����hk�Wv��H�,�8g}B+�7��ՙ�ެ������;�f����]�v�.Qn�����UY^�"C�>�C��:�:�񶋸�IG����thQ���9�qD�'}.�%�K_��h��з�L#ꐘlF��5�}�ȉ-x� ��ӻ�(��K˸��L;����)�z	Pok^�-!�%Z|��]S@/��;��ш��OiZ�d��ne�<�XN�i4��DHW^ii�C��*SDv+���`���r��{���Ȩ��>&���0�\*���J�V��w��_H�)2=e����ns��Y .����O~I�1�#�l��Z㈷t�q�J"���gt�X�
~�A���6�ͦ�)|�T�j�$���J��>usm�]��ci�E���oߜ�ƶ6pC���`L/��B����V�N
^�?�F	�,�Y�W�ǅ6'VE4q}�e0�b	�����=�?��ؿwL�Q�S�?��l�DN�'�%�h�Km(�)�m-JH�:z~�)UM�i���cM��d��`����x��:9q �#L<>���1�:X�1H;ԁ���i��[���X-g�I�&~�5Y{�}g4RV���]�|����Y�S2�B�؁C��BIy�~�E,�D��I��I'��=z��;K	\?�֔�M#�5��(��ߑ2���f:�+=�j
����^lw�9�߀���h��#wAG� h��Mi n91�#KTq��u8_�
�?;���f��Uh�'�&��F��������q2RazC����Y�R��w��gk��ԡ.B��4�/�=��'�(�F�6/�����k�6�����!���He=^-��Y:l�xBIv�餁�s�5�Wl1¹��<��{1�J�P���θ�G@��=�7C�T�=�{���nT*Hm
x��Vc ���M*����Չ!zvQ/�PX)s�b��Y��(�9�d���F������,�	�7�&f�i�OF�:����s�1�OgS��{�4�l4XlxVHYEB    3e1e     880y���c^���`�-�K����O,���sI�@��G��e�:��Kc��s���؍B�48�!�����yǢ�9�F����p�#X��O�pLq;o�e�&?I�U��n�'���ķ�sH�ȴ1>jBK��2D�	D��wڙ�qj�u	�����VҏO��J��`k������S�m  V.�.�M[%����ܼ�E���]�?��j~�Ѵ.��=:��<�*�%�QtX����.60�<��ȋ:�Q�p*�����*��g���A�6nSD�]Y< ����Z����\��Y2
��w4M�a���3�9 �LB̤Ƴ��'U<( Q�TV�>:��!1�nPN��K4X�F�g@
-�A�q��nQ]@��b%��9��R��)��]t��H��MC��N�d�3땪�X؉��5�P����z�\��`��~看Z]��ɳ|ǐ����IΒ-�q���tg�^m��Vһ}|�w���eͶ�ql������:m=0wv3���W�j����'5ng��|`��u���ldX^���@��]ݨeS�UϘ���pDB.Jڒ��r�5���>��s������Ct���+-3�����X��;���
���k ١��g}/���	�����բR2�1r�b5�+��D��`P5eᰰ��ڻ���픧�������-D�U�����������f��F-O]L�Y%uEró��BQ���j"4o���oz��,����6pbF�(u���6�&rT�o�ȡ)���L��R{��W+D~c�o
�*XCZ��sk�yO���+X����A|g�K�6�fDV���h.�8j���ۈnT��V�X fBɏ����Y���^�UP1<����*q��n+g)壗A)'�m1�*}{��WM���ʍC�,7f~�E2-�J���:��8I�s�V�OZ�d�%j���a��,k��B�IM�<hY��L��x|+�<Zǟ�m�}�  �� Ѵ�֪��̀y���ş�o���p�8���0�2�7e?�#q��~�z��qT$��]�O�������-q�k��3������P�̾�VHzo���[M���~����4ou�֮����v���G�~��Z��P��M� ��:�j0�hz�7� ��ΡR���psA1�*6_�|�ؕ�\{t0t�Y�qi;���"V��p�	�Dd�N��ǿz�m��Nsus�8+P��;�<�ݽ;s�Ml������j�" ��v��u!#��-�b���NH�����VG����&�����Is�� ޔ4����j�*���a��okj��9Q�6+[�c�Q(����ʾ��D�߈��nul�_<O�ͭ����2��p*P�*��A�ʱ�<"�M&�]���H�y;仅� � �"o+!a��9Ms�ڟ��h؏�R A��aū��¤��^�:���&k�X�L�$6�:vO�hԇy�/y��#�����}��]������[�.D3O�����鎋d?L�6��R��I��VYF���Nl�)�<��xҬ�+�-*#8D��L?V���V�s���8e%��i����T2��X���٘ݛ���,�(<!��m��d!`�9�Zi�×�d�4R%�Rq�j����/�CE���O�eqm��P{�r���׏�!4o�I��b�S�*�d�O���S{8��[���:�_[=6$B1_�H�2�}�/>K�����A�y?T�R�?-=�@�I�\���m��H~�BA���/(�M�y�d]1�BR�h�??��"F��9>p�N������'��ř"㏉.��L����b�{˘��ͭ�����l��S���{c�1���I^�X��"i�D�9�� �=�5����&.���o
"�DEք)�5a�������ֆ��:��٫�R��"������D�v�Bߖ�V5���[U��W]o�FGm�7�OB���h�x/&�����z�c�Q��W��l���#�$�{j��v;��LK|� �gZHҌ� w��%���4I\w�JWa,�.��~3K��(0��-��3���^a�]�3	�v���4RB������d��<����LE��Ȏ~ْ~�cm�!�tS,�O�\���s�`�ʶk