XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L[��Z�0�~�qN���*)��lAQo�d~��d�)��Mژm��6�xE>�d�l��M�����[��]�ٲ����:S�p4�!�^dY��-���r[>�v���*��D0�%��f蘫�Vv����X���V�<���$�-�qCtfUs֧�n?&����G���? ��OQ�pQ&� ��/�0Ą��U1U�R�2sF<���-��5�NMs,�;h��&�fF_�x�e^���u������>��C�$M�U�?��h�U�Ӝ-�]���$�(�o ���LY��txwG�J5�ļ��}��\a/L��d�zK��l��������l~��Ն��f6
]�&7P�f�봼���_S���Mɽ� f1��#T������ͺQ��-h��@�K�Tj
�$��b�K/�0�-$��rˊ�t��*5����K�QDS̨��p���v�!�Z��%����7�ku]m�L;���Ŀ�ǌ��PY��,��}�8�GO��q�0a�XX	H�Y���D"� e������y���G�P�����>�u(��6��e_ױ��N?�����6A,�ebY�����gA�0[�d�R�5G����}j:�A����C��b�B����+�#0M0��DD�����}�o���:�Y͞����5e�A ���Y����Ceג�cl¨�1ؾ�ȗ�/j���p�*ˠ��Ǩ�Y�R���T�Wƹ��,/��I. ��|+D��	G�uD�J�m�bvbp#K���XlxVHYEB    680b    1370á�k��y�q�U�|ی��E]V�Hw��,�4�$���j��ťgΊ�}H�w���
��wl0Ri�1��)W�:�_+X7�<,`�^[�B�����h�j��9N��BVRk�~E��a_$zp|R�������6��m�*?)���mG���M�ӆ.�Qu@������211�T���A�D�jq�8ޢ��j��/�ӂ͇$��	p?�~�l��"]ұ�	�"Ƒ��\�;�l�ӡ0�綇(�d�3��V��ע~@65#�"'F����M�d[I(=��f�[P�Or�o1�@|��m��ż�Pr*�Oџ!y��("�SD@Ӈc؃��"�#�;}*��]y���ͷL@G��Y�S�������k^����^oC�{��IK%C:��-��v�=�=�"ϰ���-	=:��?��6H�P�����������FzL�|j�6�g�=�-�4R�2'������+0�I���>���{["�}t����mk� ��S�U�|���	��x=�ǝ7�Ȩ��s=����r�L��������Ƴ�`�˷�mUz��e�s����;�5��踓�����4�x-�k:,L�I�H��^U�6Q��G�A�ɖ�X�s�)�U�3�݅	����	C|1'�	��v5�1y"�3�P�h-��!ޓV �v��)g���+��֭IGD8�g�T��*L@ZX�
����F�#��9�ˌI�pE�-|!e4������5� �f�����M�6t*'9iK ��ݪ ����>k2v�3T��X�#�qd����K��ֹ�^���׶o2Z �
6�{�ub��@�Jh���S×�0�r�mHީ�ƭ]J}��cw��b���ι�k���{ǲ�ބ�3v�G���Ϥ7�2cM�S#��%ua��1�]�zv���W2b3��KJM0E���Z�$�-N�gѷ����KSߕnụ�츸l5�Y�@p������B��~Өu��P�\P�.j��܏�M��KR�H������62���4�u�Z��+GD�_wCC}=v��#*	�?kq`�F�%��(���hb�wc���s���.�Әǻ�W�͗�vA~!� NbU6��F����`�����x��^��cl���4<4�+?RP�|��85B�Ko\��Z ar���-�6C�$��y�a;+n�DԨ�:ir����I��8z��T8�k2[��-�@�5��Q���j�Bő��ՙ�O|�ѓ�C82w�7-F}�ه�K�t��2�I�������Z�Ah-��F�3z�w/>��'�t�q��
��G�q���Ta�y0�	m�5QR��L�_��5�Hkk	o�^C���l3F<)&FciF���ɿ�E�q�.����k���gy�R�����<,Сol���IZ}�JݟŊ���TpZ�����Z��/���� j�Jm_�I�b�4@����m>��u��	Ə4�iB���
��[R�������H��Y��0������������<6�i�Z�vt�BȦ4p�Wy{�#-��)��(��8�tJ<(p�'��s���6�{��6�ů' 9̇���Z�`�3/���|��g���	>�j�
�� �#2GD6mM ���},�����#�]��X��J�0Ρ��9���� �Ʀ�X��?�Y�\K�N�{9��8���Ǟ VT��x���n��D���|������,(K�d����hxJ]��j��i�[�|W�<�u��[�PQ���3�� �3 �a��P��>�|G�"���7{S��~ jչ�8��]��~��� �ЗO�o�~{��;.tVIk�*���eG������*�-\����j��L� �p��7�n�����A3��"?�NDAwrـ��}+�X��]�����b\����1W�����r�)s?�DZ���'ZA,��������D �����\n����tQpϮџ�:�P�w_$�b?�EX�|L ���Lo63�;�ĺ36�0�
�§aӟ>�)S_xX��vɷ�o�L�<p� f���a�Wso�~�gO�\�zQdKJ���V�u��쀞�:�� ]w%�%��|�x?�2H_���6�('B͍[Z�~z����I�����O����pRaq�vot���I2���^|�"�o��A{٣(�9�ZUH��B�+�W���]�����wNs�,����?m0ӗ�����4;*��٫�0g<c(�/�=�ߓ>�C�*���1��D��Ɍ�C'K:M�XD�-Bo�5�R^)��3���z'���s�Nל��%���r�.h�Y��ؗ+�S?�I���?q�%:/z��^Ի��:q�v�Ƭ�������	q��|�wb���wo\:~����C`�J���
Ȉ�@.D��ᒰ.�����9V��_68ѤL�k��M��3���(�Y�9�<��;���q����wţ��:!����7��]����Y@ݤ`���0�%�����CGg��>Zh��$E,����-tH��<rK�_5ق�2ڥK]p[0���ٜ'R�BYtt�c��ө��f��o�"c~&Y���?�DI�uAG����@���n��u���O�-o\�6��$��ːI �ЃU�B�%��0��&r]�i=bN�(ԏ�)*FF�j`[S�M-�%d�m��� )K����e��vf����z�b�:v�)��KZ��!@�X�{G�Q_M��B��VZ�)vh��(��f���a�0m��g�A�Ɍ<�	�/$fJ���cY
�c�?8����Z0kp��9�@�u��t7o�VN�%t��_�x��$L{P��0큷 �z9X�H�Yٷ���t���&��Nx�[w��<�;L}�x?��v'��0��Q�$���EXX�����W��h��L�\�X�\u�аY>����ߜsFnm��+dyn'�F��qlT�?eOso�vON&U۝8P>Iۗ̕ �ᣫ`�p�y�\���o�&�qO��?�ᐛ��Mgf����<��)�2er�(k���Ldh *=�<Y�q�X��X�B��P��T��Z����n��?�|a3�G����(��v���&��F����Z?6���
V���+�V��� |��Z�_���L�4��� �it����!��F���8_]P�]��-+z��� C�DU$G�4�ݿ�:����Нk�)��Z��d�]�* "U��e@�浶�1������o��Jf���ߌ�?WM������P�����f�����z�v����2b"q��a^.ph+��9��3k=8Vw_�ʟ��ٛt�a��a�@�B�ca���V���s���Nz�Q8� IQn���eސ�j��Zf�Ҿ��'$��u�k��&��j�� �B���A�2d"�ijH�ޤ��O�Q}��ɿ5�%	�φ��g�oя�m�e3eŴ�]\`v���裣GܨQ��C5=\��!���c��O[Ӡ_�G��?Y�&M�[�C��~M�t'���vC�\��	�)��
��0-�3��;9���|9��5;$ri;������檕�t���b��n�P���~C/�[aE
�V5Ǩnڈ�M�$^�.0�4u�D���9;��I��2���m�Z��L��Dn���"=|/`�@wz=�	�L���6�v�{��K�{�	��}�k_3 �MCl��M�Ӗ/c tآ���V�`��F��]L4z���8&��t��k���sh�׹Es��Ad�"���"gOO^{<�;3�ҽ�;]�&�z�X���?��g���r�͸=���*�0�&|�E͑��@�^���䴐n�4v�E��%����G�e��"��u�m"H������,2�h���R�wMW�obб�+2���{�ă�)�ܑ��y8�b���H ��"�;���p��A2r�V�H��0U�)�H��h�0wWL;�ƾ�B���b�Y�hiuJ}nآ��}}��F�,���^B1��3HAgԹ:�A�&�=~L"�'��!*9}46�C1�y2���������r�؜�|�*�V}8'�9�mq�
�	m3XW-�e=B�8����߀��������M[$�UC}�@�W�Z�l�9�(�퍮U�0L⃧,)Y�ESá��-�ҹ��s����˹mb�ʧ����,s�a�q=���Z��<���6��#��0qi×�O�NY� Nr��zTt��Ъ��b�@�>�QV@Q�5f!��Ɣ�R��uw.Bو�."�ՙ�����E���A�����k�e����œ'��\�A$*�"������T!hT�e�ŹSa�7�\+��i��]���>	�S5"�N�w��0oo�TA0vD�9�d?J^��2�%�mV�x�v�r��1����(�M�n.n�!���)j#a�U�Q#6�#4� �눹��p����S6D�u��	���O��G䓹7��������%��TA�Da��4%��u����-_�J<"�K�5�^��ጁËW@�O�f�uw+割���ޒs;�7��a5��A�'����F��K5&��PsZ)�;��ˠ_��Ajbonmح�0�H�W��lJ���"�UƤ�4[��H��Z�ePQZL��,�ʶ��p�����\�~Q�,�ߨ:5��Ϩ��8�����	�������J;}�y�a��V[�zO���W���Cym�Q�H����-�S�C%`��g��x[M�fӢRI���lʶ��Y�a�Ġ�4Ur:�T��[�����s[��Ǔ��/�3��UZ�?��6G��o�7���P[uy��%�-aG��ݢw��{T@�'Ml�F�?f-ʛI�RrbX� P��;�����+�,$&9�%��.�A$WJ�Ɇ���#����W �<���:Y��oC�ԗ�Bv�{.��F��XYYJ�:F�ZWǼ��J-�m�l��-zd��R%��[Q�侖8������4��&Hl�ř�٬3�m1��'��#�8j