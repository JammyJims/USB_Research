XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����.A�>��-�At�<��>s?�4�N�����S��\W�����X�;bbY38�i�|�p���|.wj%ٶ�Z�
��ǠwF�:g)�;W�o����|7���%F�b�snj��F���)�=��E�щu�L?�2�ʄR̽'�M�����Gۿ��#]g~�{ͷ���J-L���hb2,�V� �خ��gL�ܢ�:Ѹ�����菦֌����(g���F~�[n|���vnQ�aV��i����0&��il���y�)��5�[B�Hk±�W�^b��3\Q����%� |7�+�;q��t�29V�#��F���눕&p������}�ڻ>�b?�R��.N����EQm�v`�7�t��Ez�W���܀�Ϝ����磌��E��eR0��5����;z����S��nS�����?�:�^m�l��(�p��t>n9:���Ol�3e(5'�A��e�ݸ!,4_?7Fpc%U�R�5�B���K9���M��a+�j�᭯	L�ruC�v�>4ї泲S�h����Mޒ����X�S��h�9����2��}y:�"�p���Z��a�@Ǆ�>��� �Lܩ������tosf������Cx�~[$��n<�����?��i���nl�����=��y�7���`�E\��$I	�D���Ik�d�)��q7s��wSP'hF���/S�	x/�[������zO��J�Fis�Gq1�������\���$4��g|���O�t?�k�G �E%Lc��`�\-�XlxVHYEB    1c52     e70�_�����r�MJ�}�k,��[Q�(����6 ���i��.wO��n<D)N��u���&������k���E^*2|���+��1����Q�{��v �qˬu�L�> �fg�u>JZ�vDSW��Mxj�!�_���`��/a�@�x�b�3��:E��ї�퓺"+�����ɇ_�A'7�
:6�-��W�U��!��H�:�����PbY|����_����Ȥ2���<�L�R���.aOi��I!�yPj�����+�a�c�I��B.($Y��a.��I`pp9���D�"`LE����S�m0Ԃ&���EZ����C0�ۯ2����/5�ʹ�X�t��NƬܬ�7&���w�A3�K�� �E��f���h�C��4P/�Q.]x� 鱯�-�,���!`+y���x�ɉ�*V�@&���z@L",�H/�)�@r_7[B���o�Br"W��2����Xa�����`K�NN��"��'�ǧ�AL{&��ܝ�Q$��_NqZw�-�U=��n+ D.�{�$}�,WW��j2�:9X�jG%v�i�����u�����f��l�	޻�
?/�/Jsӳr.V�x��b���/�/ե�ܴ��sb2`2�!W�XlA����6!�T�n���5����(���ԙ��;����q�o"	�˂�Y�i�9Q.���OM�'rȮ�/Ԩ�@���?�U�$�I�w�L�2��A7UP�>{��յx����j��_���Z�iݏ=�ĳ�d_�*Q���e3�w���㷊5� '-��y�V��	�A�۶-�c��������f1���PG=��<�?G0�����MH5��]�(��@��1*n��i�0j/Z���9Me�*�����*D	:��Ih�C���C��ar�U`��M���a2/������-y�<��S~�0�TЮlb�c�p���TSO���U��u5rw^]�CmI/?�����w_F�-���@Xt0$ϜG�~}֎��d���R�s�|	�~��#ُ�s-v���+��͌��MZT	Y��<�M�s��~/�6�ˏ���|���v~�,�2��1�����	������'�Edc�n�͡m�`n�xs]-أ�P�Fgի�ha\��I*�U�@ݘ�z��f*5���!0<�r]�)�W���F�T��pNO���'V���䶪ُ-R��/��F;�����,8��S��q�*DT^!���%qr��+��(R�Z�S�P��^j<<G˯��bH�&�\KAYܣ�n�U?G�a�u"]����A�#;�}�w�F��~�̆��y���Ħ�ՄÝ(�6�?Gw>���N������:9�_����>�X>@���X����ٵe�]�"^t�(��-�?�>�3k��Y��ĭ!����t�
>�~�ّ��CHGH����R�$���#��3�$k��4#��1��yBl����J":���h�����WE_�s�I�����v]ڴ��װ�����\���67�^K� ���yI�B�ÍH�So4�ȑ����N���bᅪ̀ ^a���g ���袰�{���V�
�h�uB�vGN��v��rb��8��S�܉�V��'������~	b�nJ�14�
[���� ���g� ��;"9"���0������hQ�G��zR�&Z�S�qS%�w�s~�K!$�\[oc����̚m�oA�y��XF:�uh`m�I�[
	tE��՚�&�B�%3�D��o�L�ʺ�z4�-�;6�b%tB?;�&���h���Z����}f!`}&O�L�T�������'��22���ީ�t��s����R/�p8̈́w����tfw�F�4��h�ht�Ω�oL�'�`�o�ek[�u�VƟ~�An\�����/��.��҇��s�h���I<,�����`��a#H�!�1�37|�զW8B�N����i+ni+�dж`��x}��&S�����.�1����m�K{�<@�Hm���G��Ni�U�|�=T��ʋB�H���H��1$m�n�!8(��8jι��;�N��/�֢�~�,�����̳.��|%*��I�_�6�Y�՗ǟ���u�K����n�l��[z=[ІTD��sPp��}��@�1ǿg�=�ngm�B^�%����M�<�Z��S��dY�:��N_Z ���� ���K3/���	��MZ ��FI�U�S/��W����5�Vlp+���$k�� �OAS�cm��MLP4!��-�>��D4�S�O�<:���A0
l��W���{t��we�4j���-;r�<&�����yb �ʶ6ü`n5�*��8�|ƏTc�;�b�cugN����-�cIM���)~ӿ;���I���g��z�<�o%�ZG�C�G��חJ��RxӨ�Uz��I��@��AS�5z�}im۵��I�yR�?�*'0d��C"���J�xD��Д3��:;���X8�W�4l�O�V:ű� ��i�b����s�$:/��͍3�VpgeK�S��9l���S�P�n��1�$�/�����z�� ��ϼ�gk�4��~앃G�M���NCW?6"T�::�aN����SWpT]�KF��/6�<c*��Bn�?O9�w
AU��_q�Q�n��Ш�ֆ�'jRf���"1�Ȗ�d��>T���\���a��z�Y�`��a�.~pn��<�|�Ǒ1\�5�i66[���t��uC�p��/	s?"U�?��Ǵ�q��9O�ww{�h�g�g���$�b���+��B�2f=��P~����K�ֱ9�(i���x�����
�b�q3(�������2(vu�3�����2O�!4^�IU������@v@�S*�����.��b��Ӈ��1F:��/C�`m�󕩞�;��\��~�������q�<�����/X����V ��I_�e��!�w�ZI�u���/���J]clv$��)�H��^�In��Ǎx�� Ѹ�ԂI��*��!(�z��M�\1��s8z�0o�v�����7��F�՗.6*%,��v"�7*��'�'���o��}����k*"�?w�[=��?;���6�k��iB�1��?��x�>XB�ke֒�'!�2�
�P� �"�%���Zג��J0�WwQ��MQ�ú��!z\i�b\�K^yZN9���x��N2	a \���ɽ�L�æ��<T�~Y#`��Hlf�T(�(�n�M:��:{˻ ��.,s�:���N&Q"�m���Y4q�m�/�
q;�r���L��/(���Bh�}c�L1��J�D@����k�:,�C�O �����{*��D��~�l���N��B���d����}G:��Ǻ�ZTt���?�����ؐ��-7���>��2��z���3z7�$j@
��ٲ����r�®��<����Lҍ��=��~8 *��w�K)U�&��\�ɧ��C��s�6$�4�3��l�G,r�ރDl�o�����%I���ݓ���3e����cƉcz�[��p��k��$$'�IlY�w�7RD��5���:[��і�S��0Yï����l�m���?I�n>x���I^��2Qž[�p�L��<��U�~�c��F�03�V�)yD��&꒙=�H�y
]j��w
��3�=��]+�