XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���	S��A��5�ƫC����5�_M��
��vi���%�1��αމ�_�5��{���5mj{�(�*@��Z�;�<�3�$T0�KFN�T�яr���a*��'���*�8��M1�=�!��e��x�~ҳ�zO�sZ���y��=�� @ٞ�x[�����zʅ#&�L#[��ZI�-lë�T�^0���^�3&�(+ܜ�r�Sž~�5}���4 ��2��rf�id�	g�uz��R��>x�=�>�'��t�g���v��`��ƨ{>�|?���Zy�߃�� 8�ϲM$[o��rTw-&���-��;z=Mi��;�Mq���y�He�*�%���K�a)2:��+��IЊ~5�f>7X|��¿c� l�iY�i��̀�c��	%����եR��\��j�R�U7�U���d$aލ�2�j���w ��(?ɟ8}l��9�p2<�t�~aτ7b���0UQ=A���{a�s�校��3W������5�5[!o�\eS���_�o,�C�S8�ǗiYi���~��3�[on��������}t��R��3��g"B���v�RG��+>��e�+���?�2��3Z�%��p�	Ƚ#�t�h�� ���cZ]g̀sJ,��L�P>���"�FJ��������ȇcȗSh"[Ч�t��9��!U��!X<�#��x��+*f�i���gIJ<mW���NO1��ai!�`��^h�\�h����	R��,�}�Q���I���cNF�"c�ђ�]XlxVHYEB    6365    13d0:G�ו���b��O����qƞJƐ����٪�j8�[�Ia5���$B+�S����r�%��پC�aK��nl��7�@�7�8���	�o˲�'��{	��xY��|	�EM_U����=2@�I��P�ja+W�!(��<\=>:��oE,G��GqW|�|*���̔'�!��z1o�E^�O%��_K?�5��\~<��i�.C"��z�N�-�U9�����}T�|1�^����8f��T�
��1�H����0�M��z����R�WZW���낹���4v�=@��\�>l��u۟�d��_�ﾌ�}Ͻ�L�$��,/"�G�ȗ���(Cni�VA��p�MR�J�����!�)�W7��*��:�r��[OL�N�M�T�DO�!���p��S�wq�M��P��&�4���i�[H�pή�����S��ڍ�_�
�F?�F��F�y����H����9vh�ru�y����dm0�%�ar����Å�����Q*�܏�H/�+Õt��/��ng�EMu쳏��}k~��J�_oХ481.���\@�1֞$�� �������t�*�!I���^�q\jYb��\x$�>D�*"�v���"j]y�Tmާ�KҚjo!%���W]@t�`�U�_֢�i	9�v�5%��.�mv�5�O�����,��Bٌ��5�qge�H����B�	�i;����&j�%�G�>(�yv)a-�����RE4�M0�[��׍�b��?o��������u(<v����WP�É��ȡ"pP�8+�y��;E+1_>}�t���kb[���SOM�"�o�щ�]�0�:%zua��R \��~v �T���	��d�z��Dk��$k�����i�[>�^C�
r�fe��H�(�<A>\��<Lg��$^Ѧ�_fǑ��$a1�Z��kC"L�j��gL�_�\=��f�-){uJ���r cM,J��gzH�2K%��z��s}�STَХs�抚Y���$�:IE�~����r���p�j���A�Fx*��0L�K�H��R%�˟��"np�-,�̷��6�<������b����;�1]�6Re9�Od.]+����1�J� �N2�K�:��0�r��-���� �@2*���y�w�nz�Wϭ�L�v,�ݿ�h
��*b
���KO�0�#��}�=*\w;-Qbk�a�e�������-�(��ZH5~n��J:}�{� á��|\`�i[�l��0(�6&k� 0̐n���X�މ�Opl2�h��9tJ�K׊�6�
����'i`V�GUT���vz� �y��O�;�F�(x�K�4�`L9�I��I��G*R�n�� �`�?�q�@�W��b�����5�x��b~f)C RX���?��������'<��-�+U����<~�L��y Z���?���.6���f��Ց_������39.D�X�u�,�u���5P֣�>LQ�I0/�*{�M��,9�si�מ��].`h>��������Y����|y�G�h���ñ����p��#H!��W���ԝ��e�a7��I�.�J�Ǆ������H�x $���*E�_�C�Y�X�K6���K��\�m��8V�A� ��_�Z��?M�ÿӹ@��8z+�s�q���X���mlC��^˺�بI���a��	k���I
U|]�|h��S�T.E?�	0t��vV���ľ���2c��_ e ���Ӽ��5@�����%��j5���1/m.f5W�#ބ�|�~52f��=_��$N:~H&��,n�>̫kUaY�'�5�_�W��Z݇��:F�rW��ֽK�P�)���]>{�&&��G���hl�0�@����oEƑ�F�Q����d?\0�p�d���aq��xO*b�ak=˪g���sf{ďO���mi��r�\uJH)2C,�>F~��Қ�X	Msg"���Z��	o�`���$��6� ^S�ޚ����c.�u��h��hpa���'�l��D�w�#�޷:^k�:��\m�"��W!�&/�g׆æH���@HM�(���R�N����]��=�">"��+3��Ť�Wi]��n�����V+����=c�C����5��?R�/������"�
�rN��B��0���m"������m~���ƯD��h݌��ȥ~��0���	@�`kTX��=2���>�q�w�[x7_H�鄻ӂĊ,��~;d��5��Bi=�?O�Ym��:�+ߍ�#1A�q�L�����	L|��ѪҪ�"��7D|�����ϒ�9��X���)�ߒrOLW@d淾�Q�XG L_�Z�Z��Þ6F]����ٗ���'��m|$�U+-1���S�q�i*=@�v������j:�_�ڪۓw����)j%̇W�*$39��R���j�{yVK���;����iM�������%�Z����������ժ`*�#9U+�D��[�CI��JA�/!C�xVi�4�7́A��9Tg�W����M8�����?<�(
b>g�Т��E��'Qf��^w����Cu�.���6!��RY�H�\��<8en,6_��Q =X�X�ā�x�0)�U>}Yɗ�~% p����ٝ��ǳ�*��`r��s��y�����v�nL3��; p;�8�mHq�3i+������W�w���{2��1���Ď���%q�л��BЮ~��E�s�w�$�`�ܱ�Z+|_*rV�[���kg�k2z��B��#@��&��L|�߂��y�I+Il�u��ט��{Ω��%�fA{�_�J��pM����&]�$th�Ϟ�@#W���j'N�z��t(��=�l�V�O�"b;`�􋶃9����?O��ZG
0�:H�c_n�@��I#�?Tļ�pf�Ou��Z�6b��T���ֱX����+G�G��|pўج^=���]qқ�I���1��#��oÊ���S�n\RԮrTbj��}�I&$�>��%CÆE!TP�ĭ�jM�\�r'0�;Z��t偁�2i��&n��8�m�vd�ڛ��,ƀ=^w������r3�t���À�2z�~;����{���0>t��~1��qē���"��O��ƽ�U�� �c�$Aw^
H-�eҷ��#��Ɠ�J���E�+:��`��ٳ�:��W$A?��̆��7W�b㜤
q��l��E/�Y��J���o���"����oAY����4�WgG蟫�3M��m2|����J�~s�E��AS�P�6&62�nZ�.��������l>h�l������pr2"9�L�ژL�''ᒅ��m���0��e����tB�D7*�A�
���brU�K�-_+%���I]uPƢ;��� ���{��o�(�u>��!Y�.Z���Y�������h@�к£�l�j(
��>���r'�7��U����fo�	@�Ό��t�)�j[�1��6!�RP{yߥ/Q5�`��1��G뙾��`מd�$4;��)�棢a��l�J>��ˎo��b������7q��T3�����\�{�~��'9��L����g("�P~1�2���,uɀ`��0�׳�4��&Yu�2H9�T��Z��Z����:G����~�xD;Y�/�TX����&H0�	l�}Y��h�����4�����G���(b�ͩ%��g�tSI3�,��h��z)�&�%��􅰝u�Q����G���JA=�x�B�Y�a��B���#}��O�G?��*$������K�eY�r�g���<^�Z�?d�i�N�)W�x���W��χ�锫4�����X�ͳYY�L}?~;[,8����b��Kl$�(׎�1���Ҝ�)�G�9J"���=ۃ�"�T6�3\0�c�û�F_�~��"�4r��A��Q>ݨW��Jsg�����"��7QvA����~�8h�%�Nu�,�Kp<[N;(�a3{.TY��CIS�f�3Ч�"|=d&ً��⣯��ШB�����OKS�CG{e��V3B��C\rv�U�of#��9Nc{`BV���f8X:��Q�J�}<(Hi�4�$��k5�`R���]0I�"�L��;�%hc�@q�0R�\��bgA3+e&��^'�����}q���z�VG��
����;X;�T&�r�E{z�m\RLwm��G��_��J߮�������u�VCy%h�����Y����Ԝ�ڭ�k�uv�`33�?p��:&�l~_�b�t�ε���eI���&��dN�z>��&��1�/~���C�9Ǣ؍�B���Щo̐�\�؝=iI�O�z������:A|�6�����ƟL�W6S?.[3.��9���@��q-�o�7k�/i�����~�5�_1j�I����˰D��3<Q@��&?9d`$�؋o�!w�K�X��,����s�>܊ER��"r��DP����s��L����`y�u�}�,h��py`��b�.�9{w�� �)��:�x+�b�$[1�9fH��$;�]�9C�OlT:�x��p�µ�����yz��2;���zbYai��m�\s2�z�B�1�Q���&dt�'��*�%d���9>��B.��P����l=��z��''�̺>�z��)e��O�/�I*�/��@���MO���.��֪oVl�<7�?�i���L2�
�s�=����5�����Ԅƪ~Fu@���n(}�����S�DNR� s��Kp�Dbh�	�8��T�i�Z���ɇػE
M�"o�
N��b�}���o�E��k�rҼTh'�8T�b!C|�~5�������;����.��+��&��,YY�Q�kuRw��4�9�`�m�gm��HM�I�X�5����k�%o������&�����}ax��
��s��ۢ̋�С�>�����WW�^�������,��i�q���E!q̄�O��V�!0��0�ߋ8T>b�PW�e�E&��3�Rf��iĒ|����9P�����4_tA?�	mY%S