XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����P��E�
���]���!%�bAoЗ-�pkڝ�H�z����/�u���#w$���#�\��b�|�{S��9�.��5+����j9�� !���c;IG�k�� V�w2��& ��ba:� 8�݃Kx�)�7Þ��w�tj�:v��DO�\������:��ꆋ�8߻���P��5n�:�3��(u��z����Ⱥϯ�;_Jm�@�+����:5�-�d��@Bx1�V���
Œ0U���l�0ۦ"���[R�h^�L3�}Sy�Tk��AH��	 Kߴ��]�� ~�����'��WS�1�:�2P�G1UѠ��)"��\.�w>��G0�<�����N��$G�Q��5>��u�?dh��\rGU_w>����k�b�m{ٍ�%�q�YN�lѫ��m���ݥM]����$�>\��y�Ħb����*�A�&$��ˇ�6��]+�}�'?T�H�޳�lIT��3P� K��i��>=_��c����_ݻ�wj;�C�E�����N�OG��H�hzk�>XnZ,����^vG��B����ݽ��F�����lfwR�g�c��������w	�|n}��-���vT���XC��qO����aC����wxs�޲���\t��P����BĹB��,�e	'OF���
 ��!����@�9����~�����K��0�L�l��rhe�>d39y�{�R�B�s�熙JpM�q��)EƁ�lc{"<�*��1��h}�Ny�"Z@}�2XlxVHYEB    1678     8f0~:�_0e��(G"*�m&h�B��RZ�_ф����6Ț��8_;E�q���$�,4&����ʔ_a`��D�C�_a�e�����G�t�K/�O����۟�K��'�8f���~�ԇ����G
=�P~��	#Lan�T�~�t�<�����WA�6�_��˿��;P�ޤX�b�th��ZECw�cS5}1��&����d'��Ě-�<�[|��&ze�<�m4f��g�j�w��Rn�{d����C�_���AJ�n<ݬ}J5u`�9�>
�qg+�Z�3>��M��u�	33g#�,P0ދo.�����m$b2�1N8Gn���:V���N� ������f_���{��S�x�&����d��
�H�9����j9�����`{�5�����"���c30��%lz�T�."��u�n��q"c��j��#|�4 ��`+��dP٫��N�VR00���k������#y�#��#hq[~AR�E���S�r6���%���Z��@C���|F ��ռ|{���y�|�V���H�lq>˭�q�a�9���e�?}Q-w��V�ۋk{?ƪ�F���
X�u�J:�7��Rd9�&�[\�w��ou����V�\�45�Vذ�0���6���Aݞٱ(��|v�|N�.QJ�\���!wѺ�`��b�
��x�ݻ�$�+����K,TQ�6���c�W�F.!	��P���q*��h���-Ɡ�<�j�q\j��g�%�>}�PaQ5_��q]�q����n.oo�㈢9@���� N1[y�2�3 ډ�Fۣ��W��989H��AsȘľ��v �;�k4��y�E�P��?]�|L��q1'�}��5+C�Q�%J��qY��gE1Mzd�K����m�8�o�Sn=��t@��>�� �f�:U�g��-K��hf��j���Oκ�*�Sy/�����E톣*�C���F!�f�&��!o�#r��CØ��<g�)��.�!���80v����4H;��C���1��|��P�.����{��?��X�>�OK=�e�Cb�B����n"�_��D�g*��� �'ٻ��R�����
d�:4��[�b�0[K�N��E��U>�Ω��)��'ǜ� =4�]�%[H�]:� ��o��z��:�L�r�^l�@��2J�6�-;=3nO��o\05�D���/��B���-�B��B���L��3�����RYwKM Ǝ�[�k���7���8��ݖ��	��/[��G�~n�츫W���Z��^Z��Ӓ����A�1�J�:�n�|a��{ĘtT���:��3A%cD�/+csH�5'm�#�q�H�l#I5\���M�"��y͚�o-k�^�l5< A�Y���j�nU��k���0%�;~��OALDr�k�տ��k|�Cf�h|*?��8ε�J�3髉�փ/Q&���ܓ:qk���2��(��u���sÚ�{�s��k����v�!M�}	�*�,#���
�:� U#m�"ob�	�+B�7�B#���e�s� ��,vP8Z����T�6n��8ak��C{����j�_(⃜�}/�N�};i��	�}�W�rS'�H����ɟ4$#���"���'����~G�]l�i�)Q�C++�w��A�d����T0��Yz7�M^�y�ua* [Y��@U��W3��
$�j�-Uԓt�����rs���cs����� <(0��ߏ��J$�K��Ux��1�6Ya`�ZZW�{0��phm`��j/�9�w��]/8�6u���_�Qm�V���|�����(|�/N_}����@6X��XUk`�E�� ��YW.�!_䅱H��������yׯ��%�']7��v�.�vRT��Ԟ�P�\r�b��"-s�(R��JC�����y��M�YD�&��ʻF,	_?f+/-��>A��Y��MQ��P���F�lύ|���9Ԍ������+��d��7���l�Ov�}F���ƒ��?0�K���&)I��5����t���� �ĭ~�U���Cl�����=H�D����v³��̊�xù�n��|���@F�	��V�	N}���לx�]d�SiܡY��;��Ĉ�v��wT?�ӏ<s��	 lM'����ZX�'}K�%ɤL�e�����-�j�W�#ӵ��|�#�H��d��{c(�������Cd����&u䰦<���Hl�#j7Q��\̶g&��h2\�!��i����+w��t�x�pj��<)I5I|�D�b�P����M�+�