XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y��l98�9�u1���A�(l�>��ƪ��S�^݁��ޓy�������nY��#�;;��h�N@��J)o��-��`6Bl���s	'�3�	1+f3r��bG��~K���,e>_΍�//���-�1%���h2�����A�H*�͑�%�.7��~z-E�VR�_c�x�Gg�:<�]R�r��5�������P5!�l��g���zA �׸4��D��=��g���ͤ�|	�V� ����"��i�u\��>�Bc�͒Eܥ��iiv|E��]8�_p)K��I9e��v�w4��s�/JI{�BvO����%���Ӣ����E`���sG�3QexTW�� �� 7�Y����oy���U:�iV
�G�Se|1:1���N�2*љ�=��g���{&
X��?�^�8.,hK�g@,�¥�"ĕEN�r�d^�[�"F�v��@��b�+�
 ��㕎���b]��H�k0�ӳN]��z'�ʢ(��T�[_!?^G����-�L�	��׾���s�vv�p$논-7���3�9T���:��B����{��$��e�<l�^W�?�
�ܠV��VB��J�^�1ǫ�Y+����˙�(�`�ˬƒc^����
o��>i��VG�j}�X�n�2i�3��AZ���F.q�o�o�%�MHy����N���L	Rs>�\�7RN�<K�8��)�d���`a��,'#F��f^c��T޷y���IA<��\��N��KmPZ�Q����8dXlxVHYEB    4f3f    1380ٱWD��,�~m��%j���K�P4�3Y�B���{��P8����� ��Ծ��(�&a�U�q�/��$rt�[O��y�=�A�,\z�M��������(D�\l��k���~�j��~�p;x!ou�#�C̄��:l}�;ʚB׬Y��������Q��,w!�![��$1��
O��ѿ_�-��*�|��DHE�Dʧ�.p��.4iRu����t�����!ݯ*>%��XX���TU'9?ŝ2���=y�>��l_|ڧ�[�� �%�'� <��u+\}C!�6�]�{a�̳�h��cL)L�Y�u\��"������a8��!�󪏁�W/��|���{}^/��D���}Ϡ�>Q^^�^JoB��3V��!�s=�}�"�|!�,gu3s2T~��!���T!�P?��ii��q��˫�씕���a�׎���[��p/�c��
�m6����C��kW��Lu��ꕭ]�Im�C2A{��Z�
o�Q���`٩�BJ{��lO�I�X�z]��E�[N�p�,C�����Nh���q��xa����`�[�#�O	��qib�?�J�&�q]�>�S8�����jŧHS%�(����1��{�ǑE[�b��j��o7k*ݪJn���z?���w�ʶ������
1�P��|��R~�'|��	u\��)�Mz9n�x
h�F���U+I��� ;n�y�3f����xga_����;�h�ɫ�z�vf���"��O��Q�!���'�P��ƛ2��Y)�����T�Vַ�s���h��ǀs�~_+Ca.v�E�:W�Ѽ�������j./h}(�3V5ZC��ط��l����B�n��hreh�����g{m�d�ũ�nCKqq�t6��S���qș�]�DՖu�6N%�D8X.��#���5�: _5�V�v�!��-V�'�G[7V�Y�攔+?g]��s� ��/����p�4��m����:���Z]�~���H҇�Fw��f�F%�Qn������H�Z�
���0>~!�4���7a�0��Y��JO15#�p��6���Bh8�De��Ti<�kZ�r�ML�+� ��E���Lz����U�t����]6�~u��5�J�|1��i�̈��.c����|��E���KI�D�'�7�Փ�O/A��J֔��r�oYޗRY�w_0�p�`F��F���L���i@��p/j�绤#G=��M�2�]�+,+��$Ġ��i�P���LgL�@z��5�7��ܚC�9��!(��{'������!��a��D�ӂ,'��F7A*��������m׭��*��-��PN8ت�˸�������Yєb��qA�)����\%y��%���ɝ�f�k��"��]���=��y���{>��^V_����T�cE<4y @�.�t��6.�8ԖO枲�c��;&F�D��0@���a�Rw�@�p){��G��}��%ncv~���k0���"�d�gQ��
3DD��[p@� 8N�I#Ph�{���`g:
O���'�#��T�y�[��;�e����V�1nfj<�I��I��B�?0P6�b�si�2,�f���bG�}z��75��I�a��ۍ7ySr���SR�H� $���U�&(B2� �Cѵģb���J��{�x'����/x������t�U<�$!x򠔪�E��BӺ�7H���M�>��o�fD�n�j tZtG�ʒ�h�I �=�`�"��J6�H�]>&0�1LI��)��������9�ͤ�n��E�R�������%��ԟ?u�y����:�8�<� �qu?��݅�V�@@;�䄚����9=5s�Σ��򸭰I�ۜ����*hq��)�Y�7�ܛ�a���7���CW�k�Ȕc��_��~�,~�o�o?�-�0�r��3f��3�
\�g.��[�4Jå+�@��}�drѸDH��>,�tj�3`Q�A��մ�_�[��E ���s�t@QRmr����Zk��;S���hpG�����OIݾx�Q)��K�����8��=�&XRf1!O��|�$���t-�[�t:�bU�hܨr�*�C~���Ԑ�3��Ղ/6K��,]��;��~�6��u+
�/�y�X���q�Ӽ����,�;�%'N������뉢��H*״\�0��=y&VD�Y���k��73�e�oYNx6���t��@�%L��p]�c���{��Nv�U���!��g�X���F"�=�r;���w���Q�d�b�`cS֗�s�G�+e������6W������6�Ԁ���)�T&}�yzMf� ���.=}O�e��Ea�h�m+r�L17�]�IA%�r� V�w{	��̄���
9��6d{4��p��Wa�Iy9�9��[��0�5=��3|�gY+G�\�FiA��y��֔�3�'�A�HR������R�Cd2����@灐>5�D��v��( J���'��I�@����L���H���D����cq�5�ve�B���B۲�x<G��c�r�aJ���3��J�;/���<`��44��|�O>��K�Ɩc3�y����Oj�Ql4�8�� �[�V���s��%.B�4F�Wk'�{���b]���'��l�YL	ʗl��dM�q�Q�\y�{�����sN�X�,(��S_^�mTi�J�+J#wK*+M%*,�:x��e�F7�ʶD�vI���91Q�$.�KQnH�d��)y�܈LrBۅ�FG���<V�CM����zV�4Z�[˥UiD�*[��N^���gq~�\�d�Q2[Z��UQ#�;��ޛ��>��=���h]��D�����h�.5�mi�,�s����� �L���PPt��:�ȭ*Xe(�l����*����������'I�p e�c�<�d�|
<H<���e�;�p�k��L 5=��d�X�|qf��ϱm�.^�Li�~W�C��a�E+ͮ��і�S}������o���q-Ĭ
\����X)b�N3:rw��斏��g��tו�Ȇ��5!������e�d�?R<V����4�<�޽l&�#x�Q��)Dǫa��w��LB���<I�ZϿ/l~��8��(.B`�9�f�a7�b�U���>ʪ~��kM���lz�Ø@����>�˟��>�4��hM�"�a��x�}��%}���|7�w��"�.�y)U��;�_=�ݞ���竞����#��ic;�	��5�Z"I|S\��e״_o[ȋT[��Q�)0"t<�/Ê/A�/� 4e7�I*Tv�N���F�)����:LI�TɫF�jچ���������#��~5��^����S�B_&^b�i���Vs#�?���"Ҝ�]�l�c�������j�;�C��B�;UIQk� ��R�\�xb��9i�$�;r�F�JD�M��,�r���3a5������k0���f9 �zw�(�?�����
���F�N*���9~���w���{Lj��gQ�Ot���Z�H,9G�s2�(�65������L�R��#��
�[�фA(Aܝ���8<2���"�i�3ء��f�ь��O���	�d?e#9ё�=�O@������Wscl���i����Lc���N�;k��E:�)7P'�O7{:c��<<Y�`���@	_�������$�s��q�≁��?�qI�H�d���h��ץ��/��d�.�T�͸�8�qq/�X��I��>}��UL�8��nb'X��!���7����q����_��m�"��
=�}��g5.� ��d4z�{d[�:��y6j��yn�9G�0˖�jY��b_H'����M_sD�n67J�
a'p]1��/��fkKN0��|��0# _3gŋFN56Țv��Zƽ�$�!�zKR�h6�=������Y��K�$�C4q��7��UY��? a$��弔jA���S�����ғ�U�Ӳa� �S�*��L��������Y���Ԍ�\�a%��J̃p�a7�}ͧ�0����9��&�k�/�8T=�'�I�6��S���e��_ݩ��.��؈���O�R���mw,>C��uŬ�W��d�
����Q���č����:�7�Z>]-υ !���+J/|���Ô����[�A#y8Y����0���:�{b���I�ğ���d%b]�>��PR݊Жz���B��2M7��4=Z�0�-^���9�vӢ	��U8��"���";��9�1v}��\ŵ��w$F�f��=#�=o�O��Nn��Tź�?��7���áT.O�k�9��H�hW�9��(5�u���0�n��C�ޫZ-"�n#�J��x�8IGe��*;�,��
Ƈkd�Ҩʕ\11Ϳ?��p�⚻d��Lp�v�*y���2�� ,���8w(:����\<4$��s��(S��A2;�y�fEU_/fw�k�u��h��{��h��~� 47/?B�Z7ΜmqEB93M�����\��{"{J�4�G�V)�#GGמ.��KSP�7p�0$s���G���D��R��N��c�*J�r�~�,>��G�lz����gk^�\Jb
,��$�cEUU�e��P�|�ĞP`G��3�+�n)eZ������������z�ܽ�a�a�6�d�i���ϨKJ�7z@�{���<�����=�~#�Ҫw�K=+��xqҩ��&: x�_���e�Zum&=>� �M���/�+��M����B�h-K�Qصr��	����(>�#Q��!h
���w7��bGF2ƫ#��;���a.�0�<������(X�M@E� \G"��KxW���PS��rN���[�I�~�����z�.�v=��������)w�=�	`�*���t�q\(%�n����iO���Q���w ��}��]�X�=�7�_���9��㡋Z�7Ն���@|�S.����ѧE�X��K������3	}�