XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���¸Oɂ���E؝U %��B]�Jx�y\��p���t4�^�.����v]m�� #kaO�s���l/�T��Ɋ����(F���:͈ÙP���}�rJL,=�b������G�+��1g��@Q`fC�a���h��)�S�M�.��>]���1M=�"���Q���g���O|\�OJ��cM~�z�?o���[����he�_�3ɬ�M�$�^ި�:1�O�lǳ-n�Ρ��>�E>`טּƤ
2 ��ř�5��3���.9s'Q՛���ln��6,^��4�僫�m������]	�x���5�;�����EF3k�3����%���a�ĈD|׬��h�����(�{�k=a��1����Ba��i���πF�GZ*K[�g�$'����|�ܱ�>Y!{���)���{{�i��O!R���m��<��ML�|�"ޖ3��@����m�AQ�:fu���D��3���ҩ���`��R�95tZl����x�tp �oEy*���l-d��J����@�~23�����2�`Y�d��M�m��q��R�ļ��"[�x!Z'$=� 1�~؏!Ӹ�4̊��
m
ϙ'�5n	�x(����[�}]�`F��E����Q'h~�9��9|*�󱈇8_.�U��s��xo�qx��]O��J�^1b'O�6lG��,Ϳ����0L����g��64��}�$�R�S�\�����k��:�=�����r�-��N+&.7#SM"o��t��K�XlxVHYEB    b814    22f0"^[������ή�u�}_�ͮ�F�F�$���Y��R�����g��z c����ם:�]��^^�Xj��;5�����U����P�s�P�ΗjbMd'�[�Z
k[Z��R!@����`�!�|@������F��H��8� =��>o����6��_��1\D d[���eٴƬ�� 8�1�2޾it3�W�97�Y3q���6��Ft%E�ZV�vq��>����n��m��O�ghn�aa;�!���.�Q�, q*�y�����'b�����V:گo�A�Ri�M�jo7ťm��ɩ���6wh�6m�)����F=��M�3r�ҡ�%�"^���թ
P�	j�ݷ��>"E��Ɖ�Q�s��B䀭��\�2�P��{Â-W$�Py�h��Џ�\�V1�ù0������W���i-<��c�^$F']���l��bp1��V��jTL{}��S���ϡ��Mr+��>�_U�{���U��a��o�0Y�1 ��/��������/�2�l�ɘ]P@uQ.�.m~�9�~P�#"���Z��)���R��H-9D�,��GIF�[l�P�.Fϒ��W��N�[�-���o�J(�� #J�;��b�����;-	"bi��d���ۿ2���>6�H���h�2�KN�R�����'��9�B�J�����K�[0)���wr"^.�3���%��<K�q@N*�{zJ�d�{�`����-Iz*�T���9�!%�aX�mT~���Q�S#����<Z�E��U�Qu-!�D!�wP�\aj�3��X,˫@o�%4%�i�%�/�P�!r ��q2z�1�HȪL�f� ���30�<��
ܛiu���T�C�����͝���A��0�I�����NJ��v�{A�/��@O+�us"���8T ���M( '��$-�u���Ը�3��PD~ZrA���H���+<p��g 1^�#zx� �Gh�s�b���2%��&�̨����Յ9Q�����7�9|�j�uRR^����&/�3��;����������3��@A���u6x\�5Hn��X١��T���B��.HIk�8�t���(�=��r��)�hޥ�_ގ��[�lݒ�dj��m��K����\	�����o��,��-�T�F9;�~��	8���w) p�|Nj�lC��~�f f�p ��P���i;����B��V��>�� 8�Xt�a������p �����>MG`���9�\w�?�I;xU�a�@kx�/G��o�i��y��3�I{�\�g?۶���8C�?	�ͤ?���INx0�!��}���U}��&�����Y�D �C*}@fn_"�:'U>Qۼټ��^����A�ÓҾԁO�.��q�������3�y�7i�УBv��3�<Hp�
�#�i>���S.�{�3eQخ^15i�]�����c��T4F!2���!�u-V:QP�k������I*pR1�&�R�ίz�N�+�����3{Ch-$S4J�k����lZ�ck�nmW&�iV<~E�~�K�Z|�+$|���_c\���3�=C��QR1�G&��WhS���!a#
�`�F�
�c&�fe,��ܳ�Uº����&�Z�??�v}��BL���*�EYس'�\_��R}&����⧩O��~ݍ��*��U��B,��R@@�f������mo�s���tànZ �	ڶ*�������ג���8���&�b����;'h ���%V��s���s��X
���]�P���/���ř��X��C;ø�m��C�5S���=�V3��HY�}���:U�k)���.o�R���#G��!�F�C-W�D6�C�z�Ȯ�5kʗ�h&A��`~��/�@e�"Z�L�/b�ҿp�2c$�#��F�:�Q�HD\�(�/̭�Q���)�����X]�!���7��DR�}Xخ>���m{�X�>Fy���4˚�Ǳ$��'�U��I�/�8�j����S�e�ZW��?�R���q�Ǘm��D�dޠ/'�lm*5�:X�|�����t��yp�k�8D�S�t:�\��4Ȗ�)��u��������@�^�yr����F�?�i����DPt�ԗTPf46K}����R��O-Z�j�X���j�qB*F�O�;�)�u��	��k� �`٬��H�C�w��3Mnj6e`̾ Z�lz����_�@��IdM�|2�Θ�}\Z�!B��5=]�7�Ś*ڵLC<$t`�E�v����K�!��Z��IXQ�m��
Z��2	�}j`Ɣ��D8��1,&-v(Q<c����ß�a��;]}_d���׭� �6tw�m�����	�$�3�*h��h�=�w�%CıK�e�?�u	���J��R�~��ů�Ɛ+�o���?jSRtL���{K��5�3�;#��?�Չ�[��KR0�u���̋�&FP��l�\v��Œ6���Y�8�Z�'�쭨\0c�����[�����K��bh��m���d��V_�Cٲ:讀�&	~?����^�J=��~�O��O����ԏ.��ޟ_IP��r`��h|������F�%���R���J�xuXkq�����X�YjrV�8j�x՗$�7�.�77�� �KW>Y��8%-KuR{K8�g�7G��·^�;��N�K5fQ�~�`��
�9�Q)x�C�s$�٦�������<C���s�]�I� �i�D�cVF�`�]���"V�ծ�
�p�xWO�}�1���vu�H?+�q��HA0���b��BO��R�=�r[�6��z�4�Fl�歠ǯ�р��Nb
!'��2׋�8,Z���g9��ۥ�8A�e��~1�`4��/�ӱ�#f�S�@�`���OI�Tx~<�z�6�:�Tgsh���OD/)�N��=�~�,���s�bK��/y3�}̈ڍq��/�p%i��#��:5f�Zi��#�6�A�����Y������8(��0���o!����_;��K9����/o�؉9�0�l6*�z�BV��}lR˱g+�,MQ�Z�eHשN���e�*v���<j��f�>Q�_�b�<���h�
��q��𡢤����G�9�4 ��Y����y�ԉq�觐!����vεX�yB3��r�w��
[�)�	Gv����/���d���}h,v�Hs>���#(���A����BD�&i��iL�oE�e��)Feq�v��ț@6�Ҡ�5��n��w;*��	
$�w�۵R"E�t�#���A�����a�i	$T'�^�_���_h��@~�|��GY�/���G��\S��X"� ��i��ˌ�/�Y��?{������͔Ԝ�[@iH��O��q҆{�.�yDA���¥��X���d�
L��+��
�f��O�ćy�@n!iO*P�67�����n+&B
ӡ�*x�;���zE�?�bi�0�s�s o#���}q;i���rwn����F*�YB�X'�X>�����	>ر{�;�h3.A|!��р�M��=��i&��X������|�h&�.C�������9�u���I`��U��zF�T��fd�*��9LF
+�[ ��ɭ�3��OaR<e&%vG����E��)����d��B� )YwY&E��86(!��~�B�i��\FL�2'������t	0�в�l춧sPt�'v��(Rc�(�(��!o��8�	���J�W�P�Hj��s8�j�<�H5յl �@��Y�K%b�٣6��.����E{�&핝��k����k7,M�bQ�u��-g v	�"��4�3-c��:�a�#���SsE9�yZ(�~�η��TX.�0)wCcB��9��V�7�|N*�U�*rP�oa��B�ۗy����5�7����uh����j�L1S�!�w�L���2Ac�/�Q��!]��bz�z?�y���������a�?~��fD�LUwkG�!�v��F=���@�WoB��
�[&Bs?�2;&�WE�a�M��G��>�q� ���ӡ�lhI��NJSgJ��;�\�v8�yOO�U׹�av�$�
D3�N� 1��Ƃr��ήȟ�t$8�w��p7>uo�=���}�KZY�&���8�|�q�~Ĵ_���s½���y'�"WSx�	�ߝw��y���ɯs�g���6t�R����'�:.la�I���N���U� ���\M���iV�UC�sH�ʙ��?�`��C2��)�������3�Ք�ֲ� W7�驠ȝ�Iנ`�^X}�a��glC4X�I�'��� BQ�`N}T���D$Y���� �/B]�-%����,6T���̍~�A�K�h.B�79�7���l4f�u�`N%�0`�>?�
p�������j�3?�n��(NF)�ϖC��o �K��!����B��(�X��� W�"�`��O��CWi�pW�� ��hZu�	����9��%y�cj���қ"s��HӞYn�U@��3V�g���+����L#�X���23����Z��=��l����J��4�4s+���d	��Lڛ�Yy� ��N.�,��,X
В�>���kn�n&tA<����چn��`�ݶ:a�©}ˍ�ȃ���}�*�F)b�,r���ǸX���Z2}wj�Gh�����m�cm��¹�U\^##U����9�V)Y31 %wIJ��Mem)�(h{�z8 ^I-�)W@Ĝ��m#Tl����* �zV%���7.Qk�_��r�֛���S0!_�XR��xmr>����������V�S5B�z۫LU��h�7O���ؐ���D�5���б;�x ��%.���P�Y�sٻ 7B����\x���������z�����Ub\�g�e���6^$����l�ho�Q�ϰk{��g.�G0X	0����x����Q�x�Ϝz�`$aQ�z�`Vy���!�����A�2:���]"��\��S+��nB�G3Mtb��~ �=�W������[�If$lX�Mrr�8�O1�DJ11٫���?������S�A��ET��4�t�p�R�Q��p��6g��=e���.w|�i1I�5�n9e�f�Y����k-Nޏ�l�~����tʨZ��Y��7v�����y�4&�	���yy��Q˅f]�k�4Wv	���qס�"5�7���Ma'�>9�d�;��g�2����#�?K�~�}R�v���%�,뛖�e#iЗH�$�����K��dps�2���ky�<8�J1J�H�=�I�zזI=�*��8x��#�^u��{�� ������:t,�,Jl�Q$�p�k�2쫼�_��zߩ���o�+�rx���������cjk�:R��#�,.���-4b�o���2O80��H(ͼ�й���&�5�SiSR$�JZ����q�+��v�ڧ�w��/A�޲�����r}��n8`�MQJ_��W�U�^��6�8#�L|�+�E��P�D�U��"�"�|]ψ���t��军��/5Q>G��C]!�����s�.o�����ϳ�Y:rO�g�zŸ�������PN���^BXa�"
�r��㸝�;;4>rK�������ml7�>5!�'R5/�9k)?�rmَ�8��0~��q����ZU�]bK���.�=�N �E@�0l9>�+僪���3�A��AX�4��n�ŝ/y��Q'�'�>��5�=���bU�4�L��@\���#�茱V@,q�gq�嬟HM������VFֹ�4��=r�\����M��<�hf]�ob\Qm��o�.:QW��VN^g�Ⳡ� ��{�tF;��K�O����v��N8��V?��mCI_�_r/��F��(�0�|j��Y�%a�y��1n�US�u�/R�Y[o��H;�<���8�7��w!�72��d�s#�K�o#p7���KiP?.����|��h]f��J>���#�]6w�F�sdQ�\Jc��y�ɪ���+p�� GR� x<-�V�C�v�6%?T��h�D8C���`,�	&S^ݳ����YR�̻D��(����*B=��WЦ!����X��1Jt3��&>m؞Ć���I��L�	l���05���&�>�p����$����z�7��P�z�6��0V��/�O &��^�\�y^����(��l��b���f-������S���e�s��6�νt���s�����K��Á��rR�G8�ùtOP�h��$e�[KRd6u=Q+��8�$�7�OqN���;D&���>3ü�bN��3�S�����`��a�j+�Aؤ�_u`�����e��������Wb�:p�طT����.�Y�$h ����-�5���:'����_�]�5��ХO<��10���x�3baf4�uV/�[�J���uJ&|h����k�W]�v�&]�5v��ǌ���ꓫ5Ե��O��������B.���u��"aU�c�-<�r0zi�4Y�бoA�c��y,lIS�v>)��B��S��\@�'�Bz�e�5��ռS_YRX�uʗ�� q���9�؆�c�㺕I�qI(�m���]�x�AkjI���������s'�$�ɑ��B���A��Mrަri��$�V�4/"P��&�L���f��{s4bC�B%�*�iЄ���Q���z�o�@������1�Q�c~���=��#\����x_������3�M�9
�蜋�-�"إ��7U�I��=ka �1�B�02B���Y�g��gi��n��'��H%k0H(^A��]�`������F�~�\�
��HƬDQ����a�$��pj�U��Q�q����i�'��-[�G�d�Ȣu�Bo�g���_���4
`��Ld'��<�E���	|��7,:�+�������k/�6jכ��8[慴3�/�^Sٰ�(L�=I7�<֗�~�(��\������R?���!�Zz���Eol�9{��0>Έix�Ũ�R��	�ѻ�#��F�s'a7�?�K&����0{���j��J?�H�h��w	�u9�P���qγZ���4^Ӑ�XJ�>���>���c�%�������%Z�� ��Wp�gQ��{;S�Ur��B������O�r"e����+m[��ôX��hW��'v΋`���0����AD$0�t'G�Rv��&���+͸x������3K��-)E;�\�i��#� er?+�+Q'��v�C/S(�[	q.^�d�ڿv�J֙ru�E����&����J��t��l�5fg��Ոl���t�1��.{ý)7Τ'f#��<��i�$�z�ug��%^zf˛�'^�ʰ<2S�LZ�/��&~.�>��ۭ�S��J��°"��T������!6S{�K^F䬺�N��dB�_5��0 ���g�x����f�3�%��O](�ͅ*9�(�v%3�ֿ�R�ϔKC���>C��\(��z�h��{1ة �������W��K�f�p4�H}���P8����?�m������ʓ�f�
�kd��+D�(��B} �3��_���L�E�]Hɝl�0�x��&�,�Į�_l4o �����r�DJ.ؒ'_�����GPh���3cH��͍刨�Y���`Q��=�^?+Vo�<&y�dm��2��f��~Z�#U4��$LB�|2#y�^�>�]y��*�)ۚ٬������<�Z*�T��w#8aA�B��$Z�'&+�Q�,:<l����bm
6���Ϸ|��:>X���W�������ղ{��9Ya-�[Ø����_��r⤦��r���	�W����]H�(���{7dVp�ԸZ:�Hơ���#Z=�3!�U�ٶC�F��J�����F���-P@Dҹ�}6�PtW��]e��f�c��ג�I�'��Er)e����$Y$O��Vm��%<*���ج~�0�(�1?h�Qz
pu>�;66��D|D����7�ԧ�������RK$R⌔�{��xn�b�k��y�s���S�t�#!�/�k����H*�Vﳑ �mj�N�!0�^���)g~�luc�/���� ]4�]��rϸ�[����Bc̱O{i��)�5��k]�16Q	_�D����c��LҾ(�����_��oIt�2߆!g"��H�^٭Y�������)��h�Tr���������҈ac��YɈ�q�8�H�~?_��/tˋ��HUq �3K������Lmon$-oB�5Zd��5%�њ��WR�W������s�Qv$�`K�~2�j�M�{^�ϗ�����E�SE/QZ�'o�������.�� �^䌉Yh�c��"x$P;2�,6��1f��L�Cӱ�T2�E;�̓
n��Z�v��: lT��8T�OG�)x�o��،�~��/qk||j<!�J����Ԡ��Vf�Y���"�z��l]���{/���\/�\��G��q�����%��
}���1"�|C����w�*>�ޥ-�յ�6��as�D���M���*�Pz�d�b��(3i������p���U	��*�i�؆�?�� {Z|	�b�\Q4�
*r$�����8Pvz�m��Hv� 6�2n��V<a�P��Q���X W�O������5/���<='��Zh�jW;����M���y�(3Yv�����)��b��K�3,`���݉3�-QE���r��(�Y�HZ�]�1(�":�x��N�*���Ô��9�a6�p��p�`
O����e,4�/��g���ǔ�1r�'�9�����,bX)��)}��D�|�1��}�8��-��lD��A�&� ����M