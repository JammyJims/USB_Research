XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b����!?P�:�z�#�I�м=��ʫ��wәܘ���;�8�7���t�u��(���r��mf��M�i�sC��Lk�����'�j��4ߜ���Dh`���u��Z��8��,�"a�>FX�]?IS�-�a�ɢvй8J��b������6�\#���Vj�xd���ʭ�k�l�5�M�)~7$^t��)o�o���
�7o�|z��b�b�t�f�e�ꅱ8R6�{o�Ǣ����T:5����C��gg:�T���Z�� ��i�Y��8u@ɄF�pzaV+��E����N��;c��Ɇ	����b��I�ҵ�j<�i�)U�ێ�΍|4�qIy�v�!�8b�/���N��{��@��&�}�LL�V�eL�K"�����I	NSx�p�V��,U������3�±e���T
�c}Ս�t�%�6�^�48H9u�P�*���b�o��|��FqI�ĭ�9�K,���;U���ځ�.6z�P{[A�+��4B߽�U���<�i��tQ��b��ਁM�����D	�ݰ`X�"����^٘8 	_H�I�rW�M���>i.թ��W��3��f�d-����#�\D�u��Iϓ:>`�@�Xl3� WB`N}R����tg�/�,G�]�,���Qq��'�`��)]�j �e0c��.��/�;l����;m����U�_/C��A��j��~�lh�x����������$��_����Fhq,��|�H�����]6K�mf{���8ҝ�l�JUXlxVHYEB    5c3f    1510�rIm��o��$��Gh�V�aN#y(�mώY.�����:��3*��������P>5y�N)a�(��'�dҟ��;��Į�����:�*�|T����}�0�C�R� �%-xo�5��K�Ģ��b�i�PT̖'8 t�*pFa�CAI'�7a�N^���ٰ4%R��E�GV}�c��+���eA�kK/��*�p>��U��5�I��}�}�*p$��6³X��o�u|�^R��~��ɑ$�O�є{R+�=2=lκ����qtw��#�gL&Ka�>�v�vz��-��u�C�t��9`����X�*R8�y(yj�KX�AV�,����8��ه�oP�/;��X�r�(JQ��U��G-ڍlh����7Ԛ���Xq�+�Ω��BK�Z⮨��c���|�%I����l_S>~��QR8	#u��|<6Ȃ���{\1�<������P�L��/W�[���u���m�]�Q\by���$G��m����i�f�09�Ô����2������eN��Q���M�.ĴMw�x�*Q>Gx���)WGՏ�{{�KQacDAVi�^��«͝`�ߝ,��!&|`�o�FnH�9�������Ab�_\s�s���}�ñh$��$8�z.�W�wh���ĸE����=�@� �ȫ�I�W���npj�u�4-��9pL�iP�B�zQ��һ]��w����z`��ʤ��1�Ϥ�B|֋�%�OIl%�ι�ﾵt)����.��{�դ�~˜�v�Z��>n3�~����o����O���hHj���\h���_�7y�y$�^�=��"j�I�;}�~<�����31�k�{�g�H�(cE��R�Jx��ơ5o�<ײ�w���཮��@sS�g-��%?�b9�#�2�#�[`�İ�<�I�rQ���P�͓�4kZ�8�7�w��^otmQ{ZeK��Xh��Y����9S�F��x@���m?��I�&�8�i$�u�����0�(�>�M�3��[XX���p(7~�+��):���g�o��j^N������ʫ�Kj_/��B�ݲu\�c(S�@��q����gՀˮ_[&6��>�=��t-`U`)������_�2q���P)�(dڊf�S�b�h��Z��k�.�Ә`��`,�%�u5�~��K��}�R+9KKr(���
I��w����9�u��$70t�s�'���4��&g�K�7� |��4!�6S�!�Ss��+·�>��G����}�9�$�V�s���V�	�_�.P��g��D�pC2����E)��\�� �f��qD=�:��h�.v�[ǎ�&����Zfz��]�6֎�1+�pj���=JM��w���\[�����ױ��N1j�c�|7�[���j$��73��!�%�^���������JĻ�����ӂTm�M?���r.2�<�>�tO�T���l�����o,�	����5����r��=�.�h��m�*��B�HJ���2�..����to��[;���R�"���r��ј�r6Q2%C`Q@Dr�4 ܡ5��%ڹ�3�nRZ����Ջ�d��'��\d�9�ۆ��m~'XH�dM}�Ǐ,*����v�����JC�xJ�μ�=�ޖ��a��eB���R3$UAKY�ڣ/m�Ϧ�(�"��վ˼
�*���M��9Oq�kf 9 3�s���e�iJ�KD�tj�p�BϨaSJP���ߛ���v�.WG�bnsD^���h�����$ $_Z�툔����?��΃݅Y����ɥ��D3�6ך��n�k�H�CD����j��U)�z��g���T�CE�\Nd.�
�Y��gj�aoY��ԡ!_�Z��{�0<"�����O����v�{��"S�mF�@9��D>KHR�����&<p�IN�j�N�t��o��䝼Jo�4�4r� j�CZ���}1(���M���1
��[@���x�ANJ�jc&1(��t�y0s�1��drs���*e������X���(s��*��\���qRr�O�'��vr4eKq�w�ZU�!
�N_��fu���`45����?_�n|��0����C�y�m�CQ�R�^\�����l�����*F��g���]�2R6�S8q<����b×��8�5��6Ë�N����^TX+Z��%-���$7Z�~�e�ՠmLԇ��/lN���][ҩ��`N���LP��X��|5;�מ��3^�j� �-�3�=��gJ	���ꉆ�~Ɛmf۬w�����~�JVƀ�����y�U�4� o"��b�a�������
V�n8NZ7ec����=0������9��hD�S1�{Ǐ����]q�'A�d�L��1��/N�Fr� %��.�Fwhc<�(H���$�Q��R�p{��� �LA��We����SL�zw���wb[(!�X���k��(��[��8z4�EC^��������X�v�t��H��@@g��ȕl�t���uA����������^�yE �*�⫥s��ω�o�$%@-	�����Qf?cܓE��^���:��d�M��0��涞�)����Lc�p�J�sF�D��;��R�u:t�ˉ��ª}C �a��PЊ*<m�"��G.�5C�|��-���H����ŲQ���K�r��4��yu�c4�7�Z��F�^��m��31S{@�zx+�Vȟ(�	J{|Xuby`�K��P�a�G�>�����ΝjZ�� ��y"�s��B8�f�hs�/ˣF ?RE�T�.:�vv�	�8��u��H�G�zd�FݠR ��JU���,�*,G�c4U�˘(��ZM�������s�)1�2�.G�O�!%;��ud�۪:�!�g͋n���i��D�8��X�ѡ� �nq��2�C��
��B�~��eR��;')�c7^�u�$`=^V�V��|�����AJ$
t�����o�^Hm�۪�ң��"4"{b�p�:n�R>�'F�@��dVS\�=e;�%`K_�G����9'Z�y���)�BY���F�VԄ'��K�Sg
�4����;�D��$`��o�����h�;�����3~���?�Bߓ����vrnf��ͩ�a��Le؁i��,����R��3K���S�������2�Kc���-/�|H�V��Ҙ����7�e�4y��̎�sqZ��aY�Y����\���]����Ĝ�d}�w?��͑��P�C�S�ʔ�Z��4�5?�i7��HS�RYlCj�;9<0#H��f�<5U��k;9䫢��uy�bw����J��/��Ev�Ҡ���� U	r�;�T�Q�bj��N�>1��<���GYD��"׃z��aY/����zJ{��e>u�L�vp)�2|�>��<y�ހ��m�s�֬��-
������3�A���p��R�	��frV���m��<�
&��z�?����9��,���� ��?���/+8�1,����'��m2�7
kɅ� �%�?�j��+���\�6�/����"W(|�ܸ�m�A�)ʹW����2_eq,����`�BPwW�5aw��s~�l)������(��B�\�hsZ(>�T��	a?3���M�q�%Ooeg�Z�1Y����:���D�t�O�A�J��{�C6;�/��2ܙ߈��C
��[�,���6vf{g��А����А������d�����ù�����~�ݝ�%��ѝ�ɾ*�w�N�����g�+2��#�DTt�U���?��3J�׋v�d���)7��;8Ne*���X�D��'a{A���
�z���B�!o� j%�i]��eۧ�8���Nȉ5wM?ہU�)R�C$��a�����Ʒ�D�Ҫ��k�6���B��!5F�������+��&u[<*�)���F/{';9���ZҒ�{��D�/5�J
�v����D��,1C2W��
��c�La���j�)��^��n�_�9ݨxzE�F��'Fy;u��9�)�'��M��������K<O���>=/$�q&�|��ż�(�����}��N��o��tyX�b��5��gp���Ը����K�(N��t��e	��轡�J|[��|#��4*��q�jX��vG��E��u�!<48�
��6i�/֩v�Y�l~%�mL�h�`���?�R�k�t���P�XS�=��*Z[��h�n�33b�Ȯ��jdwE��`ws�s������?kD�?�T�%�8��X51H(0*�(���x�UJ.���u��x?�C�	j�͔��U̔{['�ւ@t�.$�a:b��ln~I/(_�"����@���R]=?��!A�����1�J�M�K�?�>�$׏i��ރ�����a�k�A�Tb�r�u
�8�����,���o����ޏ��}i�婊OBs�a)֌(�3����Z��}l[ڎ�j���~��R�7d��ښ��2Ч�� G����l���G�wP���8�}�	9�Ga*��^�R�����$_����3�NǐjL���*45�h�w�n�AzX/F��q��?x�z�J�&���\5���Ta�9������[�|���L�&�WYe�$�K8�4
!'�!��hn=:5�9/�+Z�{t��L0�
�8�jO|KR��	Z�4 ��G��K?w�η�q!bދW8x5�W�{�����
^�c����G��of��Hi�x@z�-�;J3�kē-_݋hO��r�.b��"0ş�>�ɄM����d^r��@�ě��=�Jx���	.a'������������\�_�.����D��!}��t`�+����  �e�6�&���C�����x�����\�	Xd� �\�1��\`aࣚPK/x`\��Bi��=;t⌈�^%noKm�A����v� �w{9b�eI��!��?���T���Ēl�H��f�ތ=45t�u���/;TynM<�D��%�e>R ��#V�������h�I�b.t1�P͒�+Y�nō���m0��O�^�g`��E�#g�77�E*/�3��+պ�3e�n~�p?j��
aC�&��h
�ϋ�'>Y��"f*�M�w��F^{"�Wkb�
(���_��X�*έ�<a�4b*��R��94 R~.%2E�:�m�R�W0�p��X����1c���8�eQ�`��b��̐��d�/}��{�m�(M��т�vTTc�{yn�r�Z�3�+�[�j��Ys�O��� f m���j��Ĕ�!�)Ɲ��E��{��"~���w⹎��^�f�d�;1K�^_f�q`�G����(,�Yުp�`�������5Ex܁���zr9�