XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}u�ǅ�I�m�����i�G���וs^C�-�tTV|d���*�Z�Q_��6k���\NX�	*9�C�H������kP��~���ԔW'�R� U���b�n���D>.	]�]��@!x\�-c�q��"c�E��-H���u�l�f�pNUZ�A�9�!*�.v��()�p��;�nF��žt����]�$u8���_���j����B�r�f��d 4=�
�&�OH�������N�k��V$D� Ș��}{��l����t�E�\�G�<��l�(f%ذ�|סjJ~�5a��,ug��)� 4��1���Td��o��"!�=^�����`�9�J�䩚�Ja$�� ��diDF3M��
t?N�m;F�����l��v�)��g�8a�q �MR�p,'�����}�ǈ������:�D+"2)7������+m�9����}�Bt���'��y�u`��� ���ƿaC���������I���ڇ�7�ЏA`)�	��10-��c�<�)��RHv�O�b�iM�!j��f�n藗�ع��h�syp�6�i�Ȣ����V��˔�/`vS�[Chω�/�����Nu�"�9#q\�M5�7_�GЁ�ȃ��`��\H5���GMDl���|�o4"\˃�qB�?#��_C�8��͗U#�4ʲZM[Y	K�,P������V� �g3�VŁJtL�Wz@⍧��r�榣s�!
h�z�,�N:jr�@�uP��Z�>����@��R�:sXlxVHYEB    35f6     c10��H�v�vv6B�+a�D
.F�IDx޶��]��0Soj�[�&�7j�5N��|MꮯY���P3g�H^,�����r�d<͑�ڛ�Ϯ �K2qxa�g"�oD��]0u(H)��^;�s=jT(�.zL�8��iۅZ܎`���-/�i٫4��σ���5q!�+5앰��ge�˭o��	v��1|Y��ҖH��X���ؐ��r><h�W�pز����[<\$�%8D���= ;�V��HΧ��&��5�-8P�a��fLv}��<TA8n�Z��p� ����Gb,��q"(�à��M�A�ҝΈ�T]�*�h��\3�$�Y��x';`��e��d������ ����Ղ�/IP�}�c��J��o'�Nߧ�?��&��'.nXl��U�2���T$`��h�=�f�y����pu2eZ��k����#���2�{u��.�)n�d�k�#jg^_�z/�Fi�8B뿤�¾�r��C�F�J�.Ӵ'�'��"�7F[s���k����G�^,�c:-��D�n<c����=�Q����uju'��G1���	���,M���I�qY�:��,ٕ��<�����+��?2���O�s�L�L�W*�����
��8M=���l�V�S�'k��$�}��)-���K�רC
��[1T܈U�_��3���#�2��v-������C'ȍ��4��"7�Lō��1ˤH!�)^Dضf��+=�-jdo<�b%��|�/ YY������3.��g��_ �X�q�Fn��c]a���t�0��6��͍hy��B�)S���@F���D��&x�f�o)S�} ۾����N̰� ��{jP�!�x��K��Yp1�BÀ6�@9V��� �F�����	�fⵧt�*�����Ws����О�ʩ����7_����H���9�����,���V=�gQS� �	S���ǌ4��0���N�7;<��*����%H���7-�ؔ%2ѕ=� ����RRe�����)�#���K��4Oz��;a�S;/��'�C��h3�� +eO}}�61)+��Qn�^��-
Ե�}��]�V�ٗ���?R"^[]�Eo)ǟ�@�´�V]h��gݢ@�?@���Q^�Am��~iO��������?�RWT%����~��,hOi)g���u�}��D�	��u��ę�śt�~�8?�D���9ՔK0�D(�6Y(� T�qe�m�_d�aJ>�Y:������QVE�4�s��}20b��S@��j�=�Lp�?w�w��س���p���a�HӚ��4e�YG����E�>'�5?���̤��j�W�W�;��X�	F��d��>��Ӧ�[mP0�5��U���Ă���{�G Pk���wI�ʳ����j���7��-Pس����bp+�������@���i�ގS���
.Kk�@�
��#C{���ۯ�-w�f[�F��5�xGȬ�4:{��͊%Zĳ>��Vw�#�*�����ض�{��3�ܵCT��b�YZM=�{fN^��`5�����D�J����ū� 	��US����o眪�Z&q�]���6�^8ɣ�-I�j�`ԛy�"0~��p"�D�J�z_����7at�[�DæF�&>$m� ��T�����iwT����T)>��$�����\Q3]�O,��5�;���d�s��~�C>���rL����H��X̦m���p��S�Oz��u�h�O3x�Z�H�gx�h+9���0,� kj� �m���A�2}�6�դ@b-O�s��Ss-��;
h����0�������O�i�]g��I/������9o@��g��b�H�^E���-�� ���9��B-uB�e��N�H��k@pH8H*��rޞd�B���47�PPDV���&� �udy5: �R�@{�ޜ��1)�hK�q�~�����6���HU�.�*� �.�k�N��I_� ���tǅ�"�F����
�y�����5�]���*7_��gA-y߹���N3���X0T���'\z<�b��ڀ�W����/]��fA�'6	1b�	��-��b�k��S3;���"r)�P����D�3����Te����n��'�mF$%Ԫ��|$� ���-� ���yEݠr��@��w��B�E��S�C`�|�ő��y*���h�F��d`�a�����k)����eai�Έ4���}j��@Q����'E����x ..o/pUgY
UK�0<�dD��&�/�'��$>@z�%E���%��w���6�L){z�)92Nn�,~��`���g�E��J
� ���!����Frԥ��!������.������^c�q�@cN���#;��P�B�+�� �bԛ��"M��-v�mFA|:�`7#�XX�}F{-���V4`J"(6rX:�K��]���j����Y���� �?.�0h�i��k��~v�`�C�!	�$��L{�GB��!���@;�'���OVixlg�Y�2ͅj��;�x�#���Bk����]����t��e$,=D�6�%����ls�3\v�[`�>�N���Fމ�lt:�>�"�ډ�mܖQ� Wm�Y�4�U����.t�A�:�PO����͸1{�����r����-?�Q�����D�1J&���:u��̙aX���5L�k�դS��H�o�a���'J��^V��3#tI�x��4f�9� �����B��MvT���m��'%�l"σ�����П�$>�R@$�|&��1���H�$B9�V �O�^E�`�"�X���@:�S�0/~d��џHO���q��ס����#wO����ˁ��)���4��x9��ݨD�䦨�j4�<����Z�G�T�B�H���/G� �qeJGj+���:���yA�ڵk#A��GY���uU"Y��"���X��
�����*�Qԥ Qe^?jx��Dh����Ê���Ss��b�����N�g�'�{5��"G5�