XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s0�jHA�i3����q�!��2/ǥn�f�I��1��j#u���HL�����Hw�09r֐���f�e�h����E�ڏ_�G��T�ׯ{�/3��V
cڸ溳x]��{纯YG�}����5�s� �����F��r�
�c���wl� �j3pvj -�Mj�,d�}�w�N���ɦ�ŷ��_�Xq���lS��U/7�Ȳ�\0���
��D\�-�����P(Ŀ;���M�P� �q~xre���3Ϲ���m���x���u���]�M�R���I�����^Q"J����@�J������ۉNP�D�ns�	D���k��x1l�.��c�I�{ 
b����]�)F(P�����S{5؟Rq�~�ڀ*ťwǼ�a]���ޛ�!��K�Ƃ�D�wD�07�zq�+���{�͸����m��r�t���L��@�U��e�~���q�l���:w�Ѯi��| kaxbd�IYƭ铉3^ӵT����l����)�fU[��+x9T?��b�fq��s�7�ꊜ�d,Eqn ��)T�'���E+6�����0���bJ���Ud�[m�\�Ͳ�Q�@q��X���c�Ф����$:i����mp�ZS$�Ø*;����.�� #m6:��l7��0�Pɸ�#��'�X��A.2���N�<o�Fߪ��l��K͎��p�PZ�bK��1v}�5�����L��@V�x�jK���F/tM�8,h�ƌvZҋ�z)XlxVHYEB    14cf     7a0Y:�U�yLz �$���g4���~�A�]��ؙ��AuӒK��
��4
��Y�^�Ly���my��=�����#��#�A1���2�����/Q�w��HFd�{�Kqݔ�O�!�iW1΍'���u��s	������:\�GېoY+��~��r�V$�R\���.��N����KN�	D���l�$S���C��RfO2���a��	_���4���0�����1�n�"	��-�n�a�I��7���//�[��ք���f��~�IDU�vx��#Ű��` 2M/1AC���g�����\8{w���Xkr��ݒfeZ��rd�Ϭ�4?��ȟku<vU�����Z��h�w����^J��2�5*��8��k?Q���U��BͺL��%�#�`�C��ˋ�j�r�U7��I:��Ш�����/�_�M�Nh����% q����]缵i�g��S��X�|�TO�U�T�G4��]eb�-x7� W���U��}d�m3N������Λ�<4��ar{Т}��B��;(�)�K,��Chg�-��?����?�)���ݕ>̍�	�=ܫ�<K��|�W�.�Z>��'���p��^�b@�BRX)���<���3�+�M{�٦��	%ݷmzi6.p�X��q���5Uk��;L�t_;Vj_X�O~�N��1�t�2T��AH>��"��������`����Ƶ�#�m�Ԧ��iP��TU���n��g0 ��>i5J|
�J!������6-��-�%�6%��Y�8�_	̏��@a<�t�V�;i��`�$:��a��,;��z|H�Tx~�S��I�tO=���GєU�ĕ�r�348ƛW�d_ݭvA�D%s� ��L���DqbsRh�;�*n���bcw�Oj�V�]��q*iPk��O�8���~�-Φ,Wӟ�V���B�O����-UL��g�p�b6�G`BcNt��ҜT+o:-fX�J���%p�r7M��%�,]v�
S�q��C�����r��Ђ��%d��g�F��
�w�C��ɦ��HM���I	�wn�G�j�� �9��o �y�QdX��}�xh$�SPj�� f��9�r�}��c!��8�aG�S� M#��晻(�����Y�ϸ��0|АH��,ՄFyۦ���xc�87h����0|�Ew"�Ʌ��
� �	x����й����d���R4���<���~c�#[@Vc���jE쬊m��4�>��0
�Ϣu�ﲾ5���꿉�Y��G 
��"��ׇ	,��v���*+˗��<�|��jKL�밤�?l�>I�Q,������b�N*�0����0�J�׶��t������{� ��F���:uj��P$�DHH�>W�i�>#�r��E�O��ǝ���)@����y���?�n�^�mz�������q�z�T㈄��� bP���L��Q��Q�4�PY
�z�3����8�_wB�k�;�;F�5F/{_��\ةs�8��c��U>u�(�����N����V��$������2�!�j���U�� ���vQ���UO�GzE��4���{�h�ė���r���{�Omq��aa�+��3H^�i���=QV�~�q}oÙ&�����gPF�`<�H���q�l ��~���$��Eѐ�dT�G�O��;J��]������,�+��vƎ�35O���8���ӯڪ~G�oƠJՌ�p������tUpǓ��F���mNOO�)� #]T�c�e���:���!05nQ������Z����w[(/��zf���]fz!���j���O�>w�w�앿K��g��U)���5==���@A��5���zA��G�y{����hj�N�)Fh�{�1�Lj� ;p8<��g,̺9=�c��D��pO�q�Y����+I�cΣm
�{�Ĩ�!\4