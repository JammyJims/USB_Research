XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dABݖ���3@��R��їJ�6�7������De��Z�wNُ�*�4k�4�^w���Չ{�JS�a���-_	B����q飏�X�u����>r���UF)�1��e�Q\���p�jV��Ͻ��d�"�����P~.���>B�c]}��>�H2��)���J��o�JܖFGU�Zɯ��E��J�s�<�C�'�۷�5�z�䰟����k>���WO�wi��!`����/��(7�6Mm?���0��;�  [��M��'#n�yI&�d�[Cc�+x�PdO���|�P�?���ׇ������F�F�D��:IOM���	�wfG�?b<e�)<�j��9Y��%F|�^R�0,�ۛ�9S� k8y�Uz �ƨ3���u\q�E1���q�Ֆ��m��a6��Eb��K��7����ѡ����ŋ[")��("%;I{ftoc����3[,`��y�K;�~�G��}\)b������[!��ʑ�# �Rql��2�^-h����&�9
���ɹ '�y��4%�s0�R���I��$� ��-#�k����x�@4Y��@>?�!��{���MR1��N�����"T������$i��Od�V[݃��vH"�'�[�r���%�h��;���Cp j��(���:,��f�:#`E�xӏJ1�Ca����DrC��>�sg�
��OtŌ�	�L�����i�ּ�f���8�T�8��S�G~;F�p�}/19��C��􇄆XlxVHYEB    4145    1320��e[w�������-&��)CToZ���́"Wb�&L���GBC�GЄ	W�=��+H����vJ_!1�]s�����ʶ�k.��AY����ެ�t#%*��<�:oϯ`��S!�5ܶj9�6ш-C_se^R
a�k�5R���!.�RLJ��?�nOВV}7Wɟ����hP�H5�@��8�X�i����jO/��׮�).e0�w^�^i�M$�0�-u��d@Eq�g)��ធ��ǃO)�.��m�V�)F.!d�©��Ȑ���U����U�
!��M�$�P��^w���5	/~�Sj	���8Z̹���ޞ��o,9�㥓蝫w�Gۗ��.Y��g�})"�k���7�A,g^�c�>��/�w^�}�TƲ^~b����l&�&�����`�b�rx��Mg�4g���WKi��I� �HH��W���*�������QP�KOH����F�a�C_O�pO^G�����eH�g����9rؼD�`��떴�+�]���!��TA}%�pI�L��T���^�E5�%|a)Y�j�&���0��.)$7�b��+)�=F&G*zg�\>&�jy��d#B�gZ������W~[XY���I�3Y�^�b���pd��C)zG0�A�`a�!��I�\My��4����k�|w��3����O|��5W�rM�rD}itu}�.�R���?��H�Û��bX�]��1�ykS[��l��:	�T�V[�`�T]D��p&p%cj�f��,�늒xeK�ʠS6�3��1�1H`(7�VFV�;�d��&���y�̃���A�ܹ��s#����� 1����@A�Ʃ��;[45�N�|6	p|����v�D<a�bԺ��ȋ�6��`�)�IYf�iS��f�T+a�hc�_�7�:Eu��,L�Vخ16V�k��Y�j�B�]�HC�:�7X��M�#����|�Ңwpwo�p� �m�&;�ό��N�k	���A%�?��Ѐ�E��W�������"4A��B�Zޤ����9?M��u�GX_�v"��n��kk塈#�Gюy����ې�1s�Xj���[M�<��(��gT�}��T�!Κb�;��+�v��?1��ŗF�G��{��R�OP���rW?U`�3����O���(g��:}��d��%��j������t(Kt7���VN9��L3��S��3�Cq�gz��I54M~W��OZR������E<���O%�!A:��K��0���mZ)�5��Rh�MjG���ٕ�󯸦t�η�[!$Qp� �	σ5�8�/G�P%�p@T��_dv�#B%0d�$�v�_L�Z��b�c�۩���ujk<t������?i���T�+�鑔�"��k���T~	~^�o�E�PO/I���q+�!��\IH|Cr�L�拈5킒�5D;���)}�'Ӕ�ޝ:,��Q\�/ �\�Ob�6�q�����ǘc���;5!�:$��=����g-�跮�ت�p�����L e@(�?�k�԰���ʇb��8T����2���H�#ۑ�lM��"���F",!�]Yض���=q�2�9��}����]���E�x�v|��{7�nN`���"�s����{�/3@^��Xۛ�|P>�8�պ���?������]d
h�ZE5��]]���Mp��t���Z7�[�a����E��4�|��JM]T�Ѹ;�fH������~���za|I����As?�B�8���(o���5��B�5��j����W���K\�lxõ����vK��.ʌ���������u v�(��t��$�E��y`@��9l�41�<��7!�=���m�q��ꃴ���B�_� cW�'x1y�Q�o'��t��	��H���J�W�3�������7c?&�������7���0:ܥ��F��Y�2)�5�|E��2wv�I�����0N��k^�H_H��&�T�;�S$Ųʾp�j��j#[��K�HN
�#� +�z1������JK�xZsKJ�m'!�'���Z)����.��(l���\� ��ϔ�����$`m��@~W�;�Αϒb@�$0!�/0ດ��2��l��a'�㋓�q)΢�c��Ը�˭�P���@��E�h��t����cԍS#�C���0��'w���؛����T�!��ݙq����� [� �gY@ %�̎���Ў$�H�/$f�zۋ��a0ܜ��Rg�bY���>��?��ָ���[�ܲn^ٯF�u���#D�A�0�C3g,�_ ��7��{t�f��X^8�?q�E���4�m�w4uǝ �QI�����p��N�LA��E��q�仨W$�_p҆��IF�������]�T"]8W3o�"��M����r�;�����wӰގ�%n�7XFi���r>q+�i)��,�N��C�DK=ڀ����A��]Ũ^���tl�@J@�i�I�Zݐ� [�S���U⬙1=�,4O�O�$ھ����h<8�܎!B��!�ڣ��ΤŵD��Hc\S���Zt�z �$�o����{��4��h�0�0����|6�V�=N^�/c�È9��
,k4��׻���yc�4I�����q���w)�跩�n64̉I�B�z~�AA-*g
��oa�����Ōksr"%�4)M���xHMB#u}��� 6�r�I��)�	aB�l�X9��"��Ўyծ|�ݎ��#��%_���ǒ�m\���ur#��"�3v49����۔M �Dw�Jk��x8gg~a�gd������y���{c;Wώ,IY��pW�x�3�B!\���[ɉ
.���&9s���A�����*�>�鈗�3���o{�J%CW鵲�HR�f�,�ř�S�Q
+��
o0w���Z�o#�q8(19�q�@O
#���V��]	
��P��@�C:�/Ш��M��$�D�������/~�.���t|�Ϗ�:=Z���K~� ǉ��Z	���W������c�����ӏM���Kj�K!�#k�)ݞ�aX��� �̵[Y�nP֮WC#�q�$n�1�>�:�O�Ɋ[��!�3p�"9�,�+��j��2n��6Yތ�`Z���L~"7���諔�2��ޚ���c����>>�Y�o���dEgb�d+#?r���D��l
4�4^�=����^ �~���{z���\�DU����ȁd��序�|���bGti��b���M`���L)�b��Nt>���U���r�@f�w�r`wkQ���׬�^!4���F@�`�Rz�Z��@�--�j6$*l����d*���9U��D!@�5���9r�EE�|$��= ?@�_�N�	�
�aD-���������G6u,��[��_G�̀tU��x4e���(vTM����/F���|���Bd�뿱$e��}���Y�7%.�j��]�Ur����XP�q�ҫ�Ҳ���1-�mu��?XO��t��z�P��fL�_�#��Q,(�M���X+��V�*�ةC��N�u�R&��n7�����2�Y�CL��P�=ִKUz�������#v�3ې���(�
��{ Ix�,��õc�p���T��F#��6�KG��d����+�˰�=W��,�7
��*��2��������6"
���"�S�8��Ʒ��,��E�w�v���t&|z`�,�O�*���O�m�,�F`�8ʕa�b���oO��d��^�=�����-{ս:��v

���VB��
�0ˤ���[�����v�64���G��Q��5p�$`Dt�Z��q]k��B��"����<��뫌��{^t�ִAdC��J�l���|Ԧ�>����tņ�T�f�L�{�.�V68�����4�	Ak�E��S
q�f��,������U{mmtd�pH���{NH�dW���lT�ۓ���,��QZ���[0�YPnb��%���nh$�2$�]p�bIqQ��!Bg-��W"}\��7#I�jt0�iYLP�=�9㟊?R�NP����>�NOQ���bA�r��h���q�D!`���e7�V_K<�j�G�+��1��K�e&�c���.se{^�D�i-d
�m��w�G�㧹�14zU?{���0���:�[��;I�z�V4{�'�1}q�P5q�Xͪu��}I�֟?�]Eƒ2������"Ϥ�3�M�\���l�����Q��~E��Z��\n(jY��p����C=�B����t�h�p���m��>���$\rj�UBS�s���o�b����W0��KKG6/��ԊU�D:�<�BD�vY];+����@J�c^=�g>@�ӿ��ΞAG�lB�g�P5��N^�����W_lU��
��0.����8�J��w���I"��%)g���S���v+�l~X�0�Y���q@Be��d�^y��h��ʫ���ب��y�vt��6��+|ߐ�YN���s�HxuK	���>c�Y�x=K�m���+�u� ]���������ȽiӮ��vWv�]!WM&+G#�`�G��|�U�LŸ�}��&���A�<{<dl1���!�C���\����BF-��`�5����U�
��G�9Hu~�2m���6%sp����GZ�������@_L��#��*]�re��̊��W�� ��%��#�#�Y�9F%�޷"��
��yjU�4�m���[D�S�_��6��2�X�6|l�E���T�RbFz�%o�����|@x��1�y�����=�W����`�Y��I�����!���"�-]1I&�?߰��N��15�*�[Aw_m��e������DO��s-�S�w�`h���ej�ݩ]Cvo