XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��IB��`
�A�%u�<�o,�K�(9�$2�~�<�,��F�;��tvx��r�<s����3�N��)�j���Y8�=��GN'@6�zu���]�2�,4!��[�M�H8f ��ga³�����''6?�M&�\���r�q"�ù�?��l��]�O��;�w�����R�2K�*��^��l�YꩼDH�Õ!�F�W�G������$Ý���钶�Sn@��#�+������B����}2��O!���ٱ�{9�[�[�h'��k� � �g���P�y�]��N�Bwo��_Ֆ�~D$r_�*��J83��B�	S��:�ш.�|oG�e���+ˉ,���b���E�:�)=#9��\v�(�1��� 7i.�)�[���M��p�z7U��72lu�PZs�fh��]>򉿇���n���h'ȿ��d-v�2s�Py�4�%�����YR�y�
�5���a�M{�X��i�9z��g!�JX�{��X:�%
B�$��M<)�$��qq���ʕ5P�"vsL�Ӧ���}� N3�kl$�K���zU���ɣ��Ԃ���(?q+�_�W*�/y� �����Km$됀�U�T�H���w^F:�Ѩ�ǭq�{P��#| �f��V�ߖ�f�Ѡx7] 좫_r�}�Ȋ��%���O�b�����F���6������I@�?"��Mw�vzd�;/����B��4�$�MJ^����ѭ�ŕ&���\��Xt����A(<9=�U�
q�*T�XlxVHYEB     590     1f05�1�T��3�cvi����R�8'�2u��{�X\�u\>��lLe�ʜ7��)�җ�`�G��Tџ�����J���E��xqŊ걌W>
��� _̵����1���@l�ƻ�,&x�8\���r�}�l�]LA�TS<$-S��B�V�ll�f|�6�v]]�j�O�_{ꦘqs�m؎UH�<Q���u�e%@1E��?�#�=
��j�y�^����pr=k�TcaL����Z4�8��Q�,��(��m�A���5<)�e�#�'��aE���~ʂ�Q�/^2#�`��7D�$�X��T�g \Ryx��+yo.�Iv,ZR�*�Ѩڏg+���^���ﹴj�]�%��~�}'�٘w1 �`��Nm�%N���D��c�蔼��z�9���H��+2!<h\�Fa��v+�!��J_��=j�����$t'N��Y�6��_��,(��(��My/�9` f��e�T�0l�R�����u�f@�