XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]��VQl��N��N��*�z��ʙa��`��Oρ�����~����
��4�b��N�.��#�_�B��^=�`��~�z@a�A�_ss��h_�dZ{[l	b68�Z�2:�x�uh��n�:��a�����٥h��v.u,n`������G���n6��� �����|`�d}���a��������W��wV�����
R䜻���g�k:c �y�c<=���������R���6h"��h.��h_$z	Z��n��}�^�:�\��q#vTm�%(�����d�N,7��ܣ�×�&qg_k�3n��BKE����#ݑ(9}ػ�M���׀ �����n�ήlzDm^����2.4�0��@�b5���θ�N'�B6Y�Z����:c!v%�\��)a<�7k�����Dv�����J����&WӮ w���q�{�/}{G]�A��í�Yv��Ga�3�� S½���5��O?�s��1/�!w�~+1����^�=W�O�^Q��S�SԳ�;�2U��ӕ픋��4����	��2�2���:o�@8�l���\��n�6��h��}i���ؕn%��?��P\&�E��9�aڤ�!(�gY��������ж��ʸ��CBm�р����1\�;n;��Y(����\1#@��� ���skew�6P;V�p@rT���i%ւ+����C�r��iv7.��+�
.��۴]���U�F�&p�&[^�J�ᢻ�`��_?B)�;Uvb�<Gw ��-�{L�C~̊l~0�eXlxVHYEB    156a     7a0=�5�1hv���<At�_��`3J.A��+H˭��_SVv�����sl�!zN�R���HI�xq��ҟt���ˋQ�7�ս����Z"�~-u�&3���N����E��k�^�P��ow���*V��H���M����k�����i�m�t~��w�+�-��+��1&��̸嬌�/��-Z����G���r�?g���$l	<���T��Cby
�	-����q�4:x,)��y_?��[�H]���u���������f��x���s<h���e$ ��g9����P��s�BtL\�N��_R�.���������S����D��/��EB��C��k|�y�1��	R$#^�҄��Ɣ��.��~� �
�"nPڅ���>)�.��A�ۉ�M�/�,�;�-g��>%�WێL����
	9�?����qOLs3¬w�-��|܈3Z���%B�(t[ث���)1����~ρ�����]� �'�}H������x��.����u6�sh�����Za��i��z9�tE�<*��tl�gS�;�q^�?�LA8��pp"a��f��Y�E�ڜ��Lй�[��^�	iD��Oӹx�f�Z�R*t��%VM�=�N������[�?\�-�h�(��:� ��Y�Y�Z!HѻYl.(|�" q=�IL�����|^n�}�~���u����B>�g^`�$�0o�~��K�~��pҍ��e�!W;�qs�Q
�e���)%�>S�&_�[� �"xc�X����Vжf�W@v�9"� ���ڱA-� �p� ����d���&
	�{�KS�W[(P]@q��Q��
���ٴ�Z�e��;7�B?&4n�6F�©
���<�OwV���_��nH���I��_�la��O�K�F6��x1�#R���6�B�9���``ǁ���5p�ƶ�J���}3A\���Γp�YL���O�8��9�M��,�6�i�Tk�R������D(xc|G�<�E$L��37ݻ��G�>^���FS��C��3��h���℁g{w�,/V��|QXX�kO�V���{�Po���r�|���[
<6�-(9L�3|n#T4<D���C����B/�p�=��>�p-�k���[���H���%�
�gw1��Bt�`*gr O����*^v����X�Va���(�g+�܎D�wNՏ�2�Pb��#��r+4Qf��4�K�,��σmM1Q
�M����2�o��D�`�F�}F��.W����R�,;��# Ka�'�࿏+y�3\W1��h�5$�s5�� �Et[���F��;0p(��,�4��) |�^F����r�)�2<�J�%�:�0��L�}�Oߖ���	.�!����@�� ��>���e��.a�}a˝ƭ]���~�Z޴�nSk��%�f�{�4�?�1���7�+ �#�������9ׅ��Oj�+�}ڈY�ػ��[��@�n�~H,Z���ґj2�n�&R9į�'�H�w�g �N|�p�D�Hˉ#���L���$h���ӣ��g�v�L�Oic�HI6�xzأ�����7�n!�8kת��G��� �sf���}T��	\�jF���
� �Gggc"���q���������V�Y�L�!X��b.��\�}�8�Q����]j��� ��C3Z&[�X�oU���������y�&��j�	:���sd�����0P��1�G��N�1�4�f���G�Ӵ9>��i!���zka�{��M�G����$NW���[��/��݃A6d~{��Ȧ�������T�g� �?v�vDT��w��V�lgzi�~\��G"�ɯ|}����Y��g��6�DD]r,�6V�Ad���(n�d�z���Z��S�+�����S�7_�[3q�Z�jdi.x���u�~!��8�=�
��ϵ|X�]��x�m���a