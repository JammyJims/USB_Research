XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��� �M����0�mҖS��5�j�*�.��D�&�� 
� :֦:�Zb��p�x�3� �RX΋;����	G䲴��Jc�M�ɻŏaΑm��Pަ�d:uM;��}�"|�#ǍX~R��t�+T
�y����b�{�蠞7�<�:vU����A���(��|=��F�� ��75v ��������pQ`����Qqr� -c3J3у4.kq�i��*.&'=�,�k���_�F�b�S�>�r؎����C����09 ��X#DM�puD9|���Y���	B�g)�E7b����B��|bZ���b^��6;�o|�͋��X~���Aa�'�@kI���}���7��ܭ0,�T�dӚ���O�td±xͫyz�P:��.��U�K4� �G���X⇛}s��Z<�+V�y熦���I�zx��*��"��8d(�ֲ�dSL0Z��<�oau2'��}�l(�&��=3�"��i�lD�����1�ܲ�	"ԧ��|#�8ۺ���߄|Ӱ��4�Ĉ �u���˟P%��S'��O~����z`��|l�Kv��m�f~����tc:���Hw#I�z�S��	��5!ض��ie�����Y]/)~�*�$�D�-?�y��X�T5��t�5��V��G���XA��t��d�r�]@\o}�_�:���x����˺���Z��^�˲��k-V;�UpӔڥ��:D��'x�Gm�CV�:ϭb��h����t
�2~�hݰ�~�A�Y|�cT�L	�{k�XlxVHYEB    de54    3220�����A55)���%�1~s�3?��(��o����J�LI�5��z��L���i��ws{��0����i.-���f�����!%���]�}T.��r����Z�y�mޣ�r��찄��.�
�.�`����D��}.�N_�L��0�tٓBE��������M�+�@&j�<N�-�a�B�&�7H�2oEx��z꯰�潭�&}�I��1_��Z��UC#Ev ��{� ����$�F0ơr���W������R�Ş�M0u�"�	¾r%��ֶ�0�}U �3H�O�1Ĭ���!�4=�ŦyQ����F�E�>M�e4���c,8~3��<C�.3�>�߰X]���n�د��"Ԫ\2�c����LmL/	d�C����'�u?J����E��ء�����7�ڠׁv+��(i<[#,�$M�g@��# 'm�!� H�T�+l�LL/ns_8,������u��Fo��6�:v�q�eɩ��*N���;���$��+��Z��5��z��F�2r"
��k�(s��_������w�]�Vny8Š�t9�k�)jT�:��7W��λ7��j-��r�����s�dQ�z4Xk�Ν�K�vn��T����(���ґB?����RT�8�S�U�n(�ܠ����֏; �2��fr�KF	���:�/��k����V����U���4��4���CV�o��C+���0ZA��|T�x�v������I��;�1���s3�)"o7�d�s�7t���J{׍əj(~�()��X=�7y��ѻ������ԉa�^�^t*��A��<�%�����m��GI_��@�
��M�~?7i:���Go���g׶݆U�^ÚW���	�v�O�py+��Ou�������8O�^?�#�����%ظ�vo�((�����t˩i+Eʛ�SW�D3N�����+D6*�ТK�Ÿ�z�)Ic�͍g�YB�2�J�TAE��|�$x� I��T��Ƅ�.�n����W�aW���lG��Ė�i���	D�Gl�KL]Eya��&��$N��ܖR � �m!���=�ϑ���, ��Jz�f;ű5���5QӇc�����=;6<&m�q�gAO�DK ���~y\`�GW��A��;%\9��]-�C�� "L0�ǎ����<2�"���M����@��`��5|Y��u$C%q�7������1H��?�5�!�`F��D|����@#ڎ�%R�.P�kPC"X���K�Q��m.���a���C�ph�=$(Ś�l���o�h�y*�*��4�����Ay����D|��m��2�Z��O�n�k˚��\��$0�o��.+�[0�����2�5�����H8��b��R6J1������)ВR���n�3��4
!,bG�A &�� �f:��!8F�K,T�� _�pTR.FpM���G��6��H�'<V�r�K�k��:���惕?�RP��e�Jm��<��9��Be��J�q%��S7���\g=u���B�J�"�2?�Fm>��"��7�btl:6��+賩21���q,{�,˿��-�52*7��x�/r�	a���]Pdf׋�A�S:��i�yYq�n�fw�.�\��u�>J������"�)�݈�&-��T5� >(U[����퍨�ih�xF��71���gi��A�3Л�+ab�1a��=
���������ӏ��Y*�T>�+3�h�m�.2�ĭ�Wģ��� ��ܙ�M�����심Iyy((c�������4�p��uh�?Vd �W,��uI���!�F��z�?�_e�#�7v|s�
"k�5I=�Ŏ?*8�Eb5�V��q�ax�}�W��?��K6��B�y��$6�����0LYӚ�8U�C�x�C!<����]�e��X���B�{SS��T�9[��WlC{>[^4���L1��pR$9����������e:�s��d�B���H�HwY�N*U$F�q���^���j�%�K�mة�p��҅i�n{��V�X�����
�z�c���UI��DQ�[g!���(�It�'UG��t��A?�sΐ>�Z��+�����&LM���U��HP�u�p^P>��!������s�A�sb�YAg�Q�f�ORE)�I����������5aln^|�C��ǹv
4����O�K$�0���`k]?0�}�-Ҿ<�a�}���Űs����Z(>���p�gv�IZ�X��;Dw��+��˷�P����pq�޷:���-��G��F,L;���O}N{N����ܟ�ɨ�'M۟��V�y�^�w��#��;���33�i��Ps4)��e=�
U�Aq�㿵�5�Ś�nα��GVUo��������t��D�mN���Y�33O<{���?y%�=�v�'0�(�g$}JW��,�}���8NZ}�ֿ���"l�@;;��b�k���`� J�/h�!��]9���/�g�Ъ}��Q���&�E>>�F?�e��V�z����ʡ�w�f���VZ�Ű ~TAv�0��[&�ER%�n�n;��iej�7�H��3$
����>���+�)��gu�]T��3����H�����ݾ�\f�*�[Uy� #����Y65������ci�Uɨ���,#�:��i�מw���� vJc�Hə�9 ���X����lb�Jb��3u���56�;�k��]w�A*�\'����S]:
�ʪݱ�%q�3�{�� ����]������{M���o�&����%��T$.$$�s��Rqڦ\�2���h�P)Z��V�<|����X�~�ĻA�|=��N8�m1;NА����+A�x�/��zl� ��\SY͒��$<���B3q>��V�lO���n���|�'&�Rʴ�_�X8�������݃D�n�"��K������Й#p7{{������Ɂo�����0�m�� f�h��5����3��]}�+�R��e�>Vdj�̚ft��p��C(<7�>Ŷ�6:�+�F֏�v����\���S�X�K���T�"$|IK0:����&lp�}o�c�*L��=���!:`Jd�V�K�y�7���H��;^��T/��%��fn���jt|��x�����QR|�� �.L����@���[�V^ޱ/.���n/�Bs��hA��*��n��r}�����~�;!������i`���n:�v �#��F���J��~�(�ۻ�P��������X����e����y	���!���,�O]����@Ma##����I��@ܾj��b7���ܐ\b�G^�.�)U.�2Je��)�4%���*����+��t�U�q]|��Vư���g�p�HۉjfR�/��&�s7=
뙍��8  ��W0�o9w		��ȶ[$��q*�ь�ZHEf{�@E�0�ʞ���-�*��G��n�00>h[��'�U�5��D�[��fڲ��D�#�Y�a[�$8����V��r��
]SX���Ў���a���K��p��]V��qG����:�K4�_b�њCB�k}1�L~@f7��������+��aVi��z�^���(��Л��h(�)r]�1�Im:�f`|}��*�
0�Ռ�>� �#ā�I�4�#v�|��LA�	F��?}'�r~�|��^In>GE��;+V%4B�]N �m/�f�������/FP�O6��}J�<�H�u�� ����\�S	��*��\0�O�b�\ݢe�8vC����L�)��l���2f).�Q��~�DbL�_\}|e-p��3caJ���i��o�7~ک��[�"����>��w����$�6r�5ٓj�J�$�,|S�l��;���a@W~���7K��Y8�9J���78�kՙ~��Ť�
m�F�����y_	q7ׯR�w|�[��\n#O�Uf ��l�ȧ��qܴ��7����R��@�H���9�=�0��-Tb�0$a����L�mٙ>���ş�#��$��1��d����J�	F%z����aa���!����Z�_�(�3^���c���/ˆ'Էk����%3���f���A�n^E���,.�M����z��*ř�.T�F��Sg��3_e��;U G,���4��[�"��'��?�ec����>��\��ʬ���|D��:�im|r9�N)s^����	������ژ��quJ�1_��Xİ�����Wӷ}���,磌^6Ɨ��P���;(>«��8~�c��D͘<3>���5�X���X|Ia�K�9Pxn��=�����֘J�K;b5�	����8	�+���[��m=�u�{��g�pM�O"Vi� L֟��"m��f2	J��R0��>�~�EV7� ����q�<�P.�a�s�P[�UM���a8\)s��'�V!��j���a�;�D(1���0Z�X�2��Rz��`��g�ϊ(��ó)!p>Vx٬W^�����L����]�焊nuuh �ؓ�*��5�}÷�ݑW�N.���Ɓye[�1������k����E>*�坨7��:��
A�]e��� [_����?GM2�]&H%O����ru���u�+��5�<���nt<�X���Á$ěhqm�#��OFc�2��:~+�0�E�(=���ZM�`&��H�V�3P���kĬ��_*XM�J�H�*LF"ɼ/p'Y�ä�(�f-��<���u���خ����0T�.)�s����qF�m��5������8iR�#6�+�iM˱04	���l�BR\���bfcv��!y��� 2���ͤ�l��+S�2��u /[U|�d����\����|�z�kF$��R�N��@�Z7B.�ɝ��2*w_m\X �Ŗ���/�#Y�ʁ�/��/ZΝ�VL�2Um�6�mrY�+
��Z�m´��,
��ʗ�/�u�A��X��zz�_[�l;�s��+��8qM^�(��-qb'�s�p��2wŮ��7���jS����H�m֐&�TTX��]J m��ܰ��v��A��h���P�"��.���06:�Z#�����|D�XHA6�"l���
*�K=��Q
^��3�a�Wă(0\3�}���0LW~�CP��L�#�M���4J�����m�\ؾPl��FB���A�D�>z5�2��٪�7�,�k�G����e�� 
��ub�3z��¾nc��A���%��A�-���&\�M\��0�CԴ��%�n��_�|�ԧ��Tt�Ow�ŕ�<�c���8�' bV]����Ç�(�M?1SmhD�%�9r��01�g+���qP���`��`�	�o�e��Z�5
Q,�?�	%��yH���Ex�2_��|�#�r楔�����)��k�"��XN���_|���t���{uӨ,F���=�.x�9���x	��P�~��g�z�C�<ōxEh^&��$�޴%59������/�✔���v�qdVX�D&Ε�H�����XH���K��&pNF6/kH!�Z�J����i������%2S]kޔ��K	��lKa���B$T_�@�[E�f(b6���W:�#41��G���b� �|�W�~�4������!;꜀��d0js�ڬbI�0t&�1��}����g6��C�./�|���G�3�XY%7l'U��m�l�#�	>�rO�BZ��M��Ҙ{Kf�=�����Ed�q���w�_iDϝ:��6�Q%�n�S `e�w��]G��Ot�z�о��:����51բ&b#Ƥw�û�KՆ���g�Ջ&��F���V�9�0���[L���|�A|VDp�2�=os��NU��j������[O2�M-n|�{z���~ ���1��eJ=N��Lt���{[%��H�'�B`b}�5���eT���v����˟`������H��-�&�|p�O`2-]+O����o�ʤ@	S�`SA(��b'��m�ˉ��OU9��ʑ����jH��b�I���!��(SeF��\gYc�)1Y,�1͝�lTDV������N���Nq.�W�b�dŘ �<��#+�>{��Μd�M4HJ���$� �ܾ����n�|fBW�o�����˥�a���N����Ս�_�|�ۙD~ �h�EI�_܏���*��֓<-s��u�;S&J[��վ(Vv�g�{@�OTZ���(OG��U�/C�<�&Hz�#���/�x
�#�����px�4Q�AM���rwD�j�2�6E�g����;W�$�9G�`�_�p��PA�Ճ9Tp;Ys�❸�T\�8+!$pQ^L�59�d�e���/Q�k�˽y��ۜ��(O�"�eN��E#�S�P��R��"���[�}�O�S�p��e^ÄE���8}2f�jP�%A��F@}O��������fvZ����8SKE����w�.�v":�]Z�=����Y�0�/зV[T��D��_��?:&N��8��S{6FA�Ec
�w�+\+T5�hBp��ZJ0����G]���{B���Y�U�wl}��q-t+;{t�[$.��I�}��{�?�����Ju�ŸΦҭ�	W6�K�U@��Oj�"��b��'�c��Ɇj�,D����
�X0���q��hG���\C�	��$�6r��B]Mb��	�������qg���mW��~�6zڠ�����t��4�C�V����sN�8Z��Ҙ�p��'ቩ >�Y#tD;�z��Y9�]�la!OȨ���\e����<!�d�.�i��qnw꼶��7d�ڢB�b��JR�8�A-�O��k L��YM&����gn��O^	3��]T��>bA�6��g���^�%ݫ�g$���%�=�>,Ͻ0��#�J���e	
:�l�&r��c��O�/_��0�5���}�wjs�~�0�SXqTGc�A�S���تJ��)u��R��� �X��U&�m�`8k�6�i��*�3�*�f��t��=r���<Z�;��)w��!�Q��	oZ`�4+��%��|3/nZ��&X(N�x��˚ū�L�?\M_�	V/V6��V�>9�tF|�!j\��l���ZMO�EF�a�p���v�@��k3��|�iǭ���R�H�*��j�T!��y�Ǔ��f�[K������L��!�w�_7)�d�4�^�X�L6�/��6in��0��B�A��c�
�t!�S{� 5"�8��v�~�Y���������A-<������;�3�E{���k��.A=#b�;dJ�
j)O��[埾�l�y_X�g�Y�^�+Yˢ(��j�,-}؉��q�z�J?���aꦷ�
��s5BI��V��k���=�$	��c�S�x��$Au�ȉ=��}���D-��z�_��v�%��a��439H���q�=�
!;��8�;�! n�A�\1��wS�N�������<K�`�G
(�r&�|E2��mg)b'�K�s�Cf:geHk�ұ���:��#Y��hx�pݻ(�z���_���65�KS� ���z�J�D��L;Fu<ap�ռ�@�Â
�UT�K��V��������0�m��VQ�������$�+Mؒ�kfQU��\xf|y.f��Ȏ-bd�n.���L���oM!��4ca~n�rQ�Ҽ�K4T^�%<�+)n���Y��yU�:�A��S=����у�ݗ�𧴫C��i��Ou�GAh���h����]H�'��HQ��+К{�5�Hǐ�Z���|ȀK�Yh�V����*��Ӏ�|b��oDm4u���ꜝ���������?��X��Qt���u�%����J�����?K�ש� �u��s^���[��&��a:O��`�2��?P�U^���2���f��J�Fek\J�.&�<�i�D ���?�;O�0h^��\�p^���������и�P�h�l{AU�+a�T-��0�8�bRC�ԻL:���1i�Haey��bB�X�/b�u�����o��ەq���
���A�*�ڜ|y3����^��1����B&��0Q�g��@,�ՎUy���+���!�h�h���/���l�����寃�����D���+��-�9Sݒ�=`�(���� Ĳ�,��I����'�d�ONS	;�At[�P���]�َ%�γ	5�R,ӆ)���;�q��VBa �𮋟�bD � �π}�y~�8R��I�L�{��M���8���V�{��iJ,9�ݳ
!�����@8��,B~�E	�����?n6�2{�x��ڤ#�V�c��SHl���@;��-+K�)�C��E���-��}߃{
٤jHKc�ws�����e�{5ϰ��%�CCD�)���f7g2�󦚱�&6W6�ڑi��Z�����y��<迮\%d#�q5y�ṥ��$H�u�j��E\!�1��g�Z:�	1=	�/�>a1PEU�Sa��Rx���vG���|ˈ!��I��Vⵛ��NLgW�MѮ2w�,���佚�9��sob��m��T&�&����[��=����:a�DSy<�xz�y����Ɯ�Y�"P�����/�e˷�fx��%e�|i!:o�f�R[yƖ��&Dsx�h1�����p�W�|{�Rh��ד�rfmrTR��ri��{X^[V�p�%���pԺ5�!��LD����
H�R�E�xu�T��|�%��b����:���T����5�{�i�ؿ�#�����(㺩"�	p�3|�r���6Ŵ�D��f��\o
��AG��4�-|;A?�%@���i_�D��q9χ�ݠG��]Vm�Ǚ&�r�1	E��6�A�/��;
G$)�(	�1U-N���.4�TdV7}�h��6x����=��~���&�FL�9	q�~v�
��T�G��܊���ג����eÐ���[�V�By\�u������G���K�-亻���F|���k�L�fzSI��T��Џ��w��NU� [�=)�Rɺ���Ecd�X����	���nҏ�|{�RA�a٢6(�L9Y��o�� W�Z%��m��['��8��Wղ�j�"����F�[dp��u�2�xr�($`ԓ���膪�Y@Os�L�zS$��yL׻cc�n�K��=V[��f��\h��]��h��$}�4� �܂(��44���)J!ؕ�<�䠦ũC�t��ܮ�/�fC�Ж��75��=�� _���ت�1{�F�ӯ����k�в���T�{m7t�5"^�4�^%��Z\�w �6]l��;��)
̉6Hul�lN�:�P�K]�c���y��w!ʊ��n�6NU��#i�ϺGQ9��?s.+$F�������o�̾�hX}.w��j3��g�B��4{�-OR�����ґ��}���}���̮��Ģ��q�,Z�A�d��Tm��{�8�z�\����=��zMa+t��"���S���R7����/pm���Z0S�A�ۤuT�7=C��;,%ہ�6��4��̰��Mp����m��T����T9�:@. �m�6\R�(���m�v���������Q�7��}�wǚ�Ǥ�������њᡑ�Ȧ���0 C��4�,��W�vH�(o�_��l��*�}�"��/��7�W�F&ݏ���G��TT�+e-L�/�@�AgG� �4�tgnߓW�(��s�*7�:*������?�0�tK��(��Sc- I��eb,�c�"�`�*\̦�	ۧ��LNɜ�w���qs�i�z�G�Ȋ7@��$R�M^�����Gg{|��3���q�p�׻%�yj���\u�1_JbU#3W���E�TwO&L��L���pv��x@1�^Q��Y�҅X9C�1)�-��"K46����~��:�t�֑�r�V��>|�a-m�,��w��T��֤y��-�z���h��H=�OB��5+�<��`�:��2;����ިTٷ�%@� ���&��X�|��et����D�?�p~_��x��ƛd��E*�n���ɡ�������v�Hb$�Ag��
����VWp�}c�U��O�X���D�=nd|��čX(�_o�%���Z,;Y�n-��f s�X�x OX��,��a����8_��w/.�F��\�DK����*�������XD0�����"���� ~@���0}��:�v�xS�?Ӟ�R����qe
0��E\��O�R�u��qmOİD_����g�S4����D�MLi� �B�e3��1�&"E���;2��Y�%=Xu��g�qI\C����[��R��fmX*8��+�Qxg�gS��T+�8�6t��s\�!?Q}�)���w���Ȕ��7j$طf���̥&���L^Gw���P��/��pH-��*�
��iS���$ϼ�?gղ�Dk�����a�Y~KAΑ"���.���)����b�Pl����)���4|OQD=��\q�w'����]�NοE��q�+�yn7#s�����1�F��2`� /�)B	�D����
�_0���$9�bg�!�:�tN��M�4��Ra������I/�Å]|#�%|i_þ�Je�.��29ڇ�z�#�������L���D�ZS�B�nr������e,����vaB5,���9�`����zPDO%�3��vRY}Z��������J�*'
��o�$�\�IE� ���*{��̷��o˯f����[b�OH��{�P���F�e8?Tղ���҅�t�1=`
xA�h���z�^�D ���}͓Q�f��s}�z(%ݲL��֦Y��gjI�K I�� XN*Fq�/˼�!��N��g`�� ��}L>9|~��9x)�1R�|�)��� ��M�[}i���'w�ϝCB����1����{�G��HK� �� �&cz�����=p���-�w��o���pJ'����8n���N�p��G��!a�`����V�����v��\[���d9���ҙh�n�c:O���PL�Q�Q��8�}��pJ�/� j�R�v [�ޙ,��*��6FJ�e#�L�����2ˇ�z��S#�f������I-�~jѠ�XM������ =�h׸�_�%-k��0�3�b٨
s��N�$��)��`����8S<�|	�D[�Y��|�3L%��85����r��s��ە�]�|�i,����_=�n�.[��T[�O�i�#�)p���<�MΝA��Rb�b�PP�h����s�*���2ń��ݎ�h�b�(�kG���zf ��?��@���BE�.h�{��L�C���$e���*��D��	ͻ��&�w��^����!���g��?��B�hM]~��b�R	Lp���h5�S�֊� ��<��G��R���ֈa���ƍv[�KӍ��}���$�O�}v�5#���DHl��/��8�dШ�ք���\5��c�_I'��fS��S<��
uOdsL��.�sA&��Q�2�%�P�ՙ��~A{���bxG����b��Q>�@�]!x��)�WL���V��1�(s�r��抇�K�Gt6"�(Ճ�(���Y����;�-OJ���~2L����b�yw�����3�"v=2P%x�j����Lm���*2�o���6i��}�*L ��x�
y�"�*06�ϧ���`o���f����ĥq1r��B�َN�w�X���w���L�����Q��W�xkl߂��dkCp-��1ls��ޮ�h�o&8�PѳH�Z����;��tr�h�ݐ]�$��Z>���9�b�JI�~	 ��׵���=e�9�w�씵��/q��u�Be�!��T�����롧9���$J�I�'�q�}��a����ੰqN�8Ú�ז���ʖcqa���J�k3�c�}X-4�8F�5��z��[�g3��������).�b�ޒD��N �[.,T�&����[��{�c㑺�ʷ�-P��쳔\���n@� X���}��*,-�K��i�_��
���>��W�TaA�Ned	���,�b�"�R!{�����;�:�}0�ڟ'<h #�@��Y��
����4���0�����+�_	o����������Kx�j6̂�'����7L���&�Z�9���S��Qp�u����:\nP!�'@�.��{��O�c6필���J�GoB1.�%C�`�Z��gL�nK/�J��QΡ���? �F��ւ죺���ӇNZD����p#�*��,���
���ϕ�aa����,��8�9S,ɵk�A6M�G$����h짖���(��7�F���������o����.я�t��1�����G�웊�pl������2���	r��1ԪwI�QnQ��2��r�|o V��1N���K7��\�)&���ò���1���(��pG-,l!�
������a��� ��wg�.�1��� ��!Q����8��ۧ�:[U}�z����hw�Yp�o���;$��A�'��1�="��맓��f� ��J�M��V8Ef�Չs9�?K�����3����Qʐ,X��D"�7^��֔j�'T!�$>4��T�tSV�R��	ni{^�E�htÚ����R2AH*�8�1��8���o���/������h�"C�d�_��&\2�M�a��BP�\�oS�"���axG�xX�`� ���[�3���<[�W�vg29�&-v�k�����?�[i��9��LOjj¾,d�EC�w�����