XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����UYr�"֑����q�x�B`��*�<��7�� 1{�ֆZ��RW"��iVgk>�;�C</��9a�i�7��!��s����ʝ�"�|q�R��q9�.�V%Y�S��N�@?��?�].<8py�i���(��Z�t��I�r�^q֖��~#(��iu��'5*���]3�R�u��&���D�w����_�@1A��M�Dj�4&�<�����/Q؋s��V���J��9م�Of��������sڂ�Sq=L@S�G�6�%g���J��*o�K��aHt�Y=|M=����_�6>$R�%qb���tf܏�����;��;�{�D����u��d�|)�4}0���ɵ2VWn2"��:�(�s�k����zψ`�Oko�D��&������GK�����i*{���S�}A8�W}�Y���dY��_��K&g琓B�����t�H���Uu�&mK8=��À��d4-6hh-9v�с�p۶Ti��.�r|Oj���<֧H�Z�j��c�o�"I�`�TNn���D�ʄ[����彪`�z��3���0�|��� �ൻ���9�bU�	i�F��"Y��nu��2�D���a��Lr�kb4R���|�p}�[����v\�h�Y����-$4����G��.8�$`��Uv�H�3͋�?��!�l4���c�=+Ծ��d7 ��!��,^"��S�3�N-��M*ɚ[t���.P��Y؆f>�R���g}�lDXlxVHYEB    10c4     690���
���6����^��V�Zc�n%4.t��KL�f�W�xiC�N���kj��K:q^�JO�&�v�{���ގ�E�6���>��&��כ��6Av��;%]���U+s�ّv�r�I�zN�D쎦b�kQѮ��M�$&��Лc�l�����{n���ԟu�	T��O���a{�l��z�[�����:!$��9��6�	lI��N	����F�}Ya�<���Xy����}��,�:.:?y�N9J� �;f�)@����y��'��֢6�Y�lᅆ�L�`�+��<� ��I����O:�h�P�x}(��&{aV���@0_
�k��UO@�y�h{b�Z泇�7rq��Q@.���'�Sjqg�)�x�0@��-�xhX�]�C��7�^X�M����nA��Sv^Z]*�O�T�v��(:���� ~�m���� IW��Z�t�e�w~�������"�#��[h���P]��"��;(�b�90��?0:Gў��'�����*y�V�=�/�.�\�	�T|6�^�N�E3E(��v��1�"vϣ3���\���ն�����fA�r�*��9�$���>�0�~�����@ǳ�7B�2mC���L����Ap�<2\��4� ل�&Sux�/u���7�h�}>��R���LL_���c��ڒ̵�t-�2�8����q��|8+���
��q����f�v=H�ƹv���b)U���h�l��r
�h��="����AhxRj����7Ff�o>�R��3+�|�x,�E�Ȫ�n�p��a�q�kU���LX3��$�I�}&B��9�]��S�+;y/�EǻCh'Q�כ���zW4��m��WA�m��q@�Y�v���MM*3��_݅6�o`����#�ܰf��q�����A����aiw�Xv�����_�T��ͳ��s�
�K�͑����~�b�P�����l bӆ�<�wuލ�@y�ә܌Gs�M�>[ǌl��EL�	)i�cU���C��G-_���u���1�F2�:d�Ҡ߲��	�݈��ET9�ل:�
y¬��,��ݐ<���}��_vȄ����6�\��W��> ���5��2gVH�Ǟy������2K�^���JӀQ��_�FP6:�]Pz��0�e�a`25�p��9��̒̽fP嚛�t[����<����#��$Iys����|+;�\����q��x��v$2�B�r,2�J�l�~ϗ��=['(+�uJ[4�F�c����wr㬙��#K���ͥ��׈�݌�q��`�t�q;�@�=>�����a�'J���<A��R�@����tݪ�9V�=�7L��0���P<&%s9��ȱA�D���s���{��ް�ĿmY~�ʪ��q���S�7Z�����V�(�W�	@o�B�u؜�k��	����sQm���(�d~<���0�`���o���|�Cʝ�l�{�<��Ҏ��ѹ��r�zh�Xj�-G�S懽*������h�捁�����LH���mU��Ѽ2�j�w8�Rz�Gbƭ�m�A�L6r�Ac���p%O}ބ	�U:U�~����0eZ�<����&�t^4�y[؞$~E��lI���8~#�ou�y���~�L*�d{0݂RBD�'B[��-B��y-U�u",@