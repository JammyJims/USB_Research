XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����T��^����@%B��u}���f~D|?��Q���ע] �o�^�Iz,��v�n�����wz~�<SF���oY��@a�˷�N_���!m� ���p���F�m5�c'���T�(3�ȇ��)�]Y�HSE��V𡸦Y"���$���x}�m1�S�D_%[y[-�պjt�cB�&�bbϠ=S駄C`Kf��xiβ���I1pR4p]�7ȏr���j(O��?ʃ�Y�*h����u#UZ�tӫݯ���P�P�]�?s��Ҕ���B,�V>@B�.����u��-i�5� :·�1�J��h�[\$��w�+.)�T;Å�2+N$�޳I,��=��X��%��b��[��K�,��p��}�zH_�����p��rγmc�i�fn�اM���]��s~{s����%�&�H��t�/t�*\:�k�S�״�l/�0�w+iy7��L���o��5��	����I�>�^��(���&w�+�o2rP�{�5�Y���Y�sp�RNq�5���f�&��
;kQ��{�`(C��(�?���^��K!sOtFDA����w�,�#�8��i��cɰ-�$ >�؜��U髭.6��vɥ�>����ػ�{��v�n#��Y;�a_ɘa��T��&��@����}<��f��[�>q(]��<O��>��_�El��E���ICo��MH���j	�8�4��@��|����iv�+�����Z�I`�
��E�4�K]�M���PL�2y9nd������L��1>��Z�u1�M3XlxVHYEB    32b7     e90�7���.o�&���m�bZ��aVˏ\�����-K��I`(��T�����p�"&� �l�u�1���8������)����q-�l���3����54���+��qݑ�s���={ҒV�";�%��*4T�I��R��3s���J'��&�����8�cA�/`����l�$b;2��# (�y#�]-јD�/I��ڈ�b�m��Ь�N�����+Yp]=���9� �U�{�X�b�q��|�J�0�:�����XJ�FYt���Aג�����E�]���l1�S�2�~_�4c9�tpK��c8���:$:����2�9> ����cfh��!l	����8��穻j*m>��Dh
x�*^�)bw��t;�BG�~�o��"��;�O��6:��
�+X�؇WFz��,�t��;��Zzk�\�;�Ө���X����D�%�r�mK���d����n�����Ǚ�[������B��}U�EJ�3�}��ܱ�G��	'�9xϠ���4�D��W����m�6������n���?��:�Z��@9�#�ݤ�֘�/1O��U$Q�%���ᓷ�[���pq{>�,(�����bv�%�n�����8Q82�e�7��p���
׾!��`Ҝ,�
z�/�1��+��+|��i���qX2��}���j5�{�X��2�bX��	L�]��	��������"�9�0���e�HM��	u��� �`P�D)��� �Q/) ������9pbz�u�m�4����I� z��$�ZR@p'<��y� ����@_��50��m'�)��B�k��*\��݋c>^L{O,(VT|3RE��k�pc����x���5�O��X�>�ƨS����^���$��,�	l �%��Da�bI2E��tֲ��)�|>�
��TZ����xY���T�ą�)���Y��ql)_
v�ukY[��r�/ā��*+r�2B� l�n���(_Θ�{��Q��ǁy�\�en���h�T��-�����	���@�*U	sld J@Z�����(>�������-gg���Xч�я���}B�ĝ:�=Ca f��$_2<��D��=64��ۙύ�ӆ�0��dcZZAtlC�&ϑ.�_g��ı��r�`�[�F!,	ƀۢ����*�2�� �~)p)�:M�<� /�6�s����	#�����S��x�
VN�(�Ne	t�cӯ�2�L.x2,��EQ�d���N�|`zc�j�v�<���io杁lʕf�<X
���Fa�c��Co���vL��-�u�=]����0�}�:��t�%����1Y�ۂC\`}.{�׈��@Lo���j��{�L�����K�m_i���jKD�m�C�q'�k( �/mq�G��C�ht$y�z�2��4S���U�?�6pWf���Na�#F��.h#�ˍo>��\*�̓�j���cBJ~�N�xF�I�ϗ��0 �Z�y]j� 6�1�� Ƭ��c�7s��yb7oP��M�?�4$%^ʘ"2z�"�@�h���6�^Q��"�g{�5>B� A�4
��K%e��W���md���ɬ��-�|�\���[���*�<��6DM�L����&��Wdq��Y�C�.���8�-b4��-A���R��B��\#*w��2٢�`k&�_~�$��O������A]���}b�^��M]�s�2K)_P���rI��T�j��5�st���op�����t�c�=�����ȓY�Y�3�B�<7�Tf��F�K����k��e�I��f��8�0��T�*[�O?�[|`O #u@saATq���ª_о��b���[��c���%jg,�%:�o��4�h�8���zq��u;��(w�xW�W!�P,'n�QPJ�_�}��"�yUq��gw{����4J��PƕtH]P��2��a���Z��g�2��,�A�l���A+�@�o�SglWe��Ƒ�<s��(�..����:�&�}Xe�_�<���1.aoy�p�{���/�ސ�!K&�����DB>�㺦�Ț�D�K�*����I�n����˽�_�S(5 ����ci��:A��;�X�G�jCP�]��vp�5*�U����,��o��d��G��G�D`T���hi�餣��b-d7��y��ۗL���To��7��Q8�� Ԑ3nl�b���lXd���F��H���G�9���/*��1E�Q�e3v���&���=cX,����`�$���!QB��=���|�T���kڇ���=�]F3Li/��W��$����-�Zz��ͦ�2��U��1l>��F���>�H�F�puK�P5G ��,h��E�{:��@9��+J���¬��l�q�u�)��)˕,�1dZ����d�� ���'hn�K�3}�o\^���T���g��X���?$0��	+�:|ѧ.z�L|[�H��
x�cg�ϝ�6�SG�v��p���Q��Ѳ>��^�I�9h�X�nMB��6����&%����x13��W��CK�Xg�/I�6��z'u�+�El;�?H�~��+�$�Y��$]��_riR>$=���|U:�.{�*�ҶH�X��G�(�v�'f@0���7��{v�'���I]��؍�q�� �3�_�WJ��. ���mj�Mn_Q��Yr�G����UW6I��i4]�P���M=x�q�F[E��\L��`���NB]�׀o��y�N���e}v�jrxccriڵfO�1_��>�T�&�B�i��q��v^���~IF�r��m�F8�Oj��Tʋ=�^��E��CD�2:	D�����L��E���:��)�j:��db�r��v�(FuG�к^A�[���r���ٸi��ߓ���d�~닞a��ڋ	�iiO A��wE��)�Ҿ����7�s{�O�3�v�w'������ڴ���tz!)}PN��3&%�O�a^��Nv�(кj�`G�ݱ(�ш�r�GE4��y�#&R�L���-£�ʑ�������`�n~������RI���'D���^�-������ (�nU�S��;	z�V+T 8��� hh��29L�I"\dN�N]�y[�$#/��[_��K�_��M6����~���>X��5W�$�B�a��Cb���"�����Y���+O:E��Z'��>6Rw�T~=cY'=,X�!�ȼ���{]k��s5`�KRfP�����<���	� g����&jp_��:�RN�;	�Z��RI�����Gq4r�w$؎�K���g��2�R�gc�H,�f�"�k7n�����n+�"��	�J!��i�4By[ih�)[ �wڊ�8���r$.R���69!��v�Of)�*IЌ�K�oy)7��wc}���CM/�ع{m�<K_@_�Όʛ�I�z �Į����L�"��a%m���-Z%*;R�����<��Ag����Wv��Hղ�1���\�|?D�e�"[�@]��[#�o�VvIf�45'� R8����O(�d�`�b���1끣spS(�ˢa�<G0I�&�6�;���삆�FmOI�%���R<�闢�/�/��U2�ю���N�G��Y�`��-�k�>��4JR_���p�-�}{���������{��	�.�;r T� �U�c�_�] J�:�Ma��-�Z�vږ�*w���4ȴH3�<�VS����)F�