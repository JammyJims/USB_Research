XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���EntZ�T� ֆ�o0Qa{��X#l��dr@6�j:���=l�mCm�_���fo��h��vf��qb;뤬51&x)�XЈ/������$���cw��y�/l�鬠F_��� ��Է�gq/�=�(�7~���RL��"�M.�ݹ��}���*����;�U�"�I�-��F��¥��D��$�a�G����d���|�����Mjv_����>�{o��>xi��-���G���t��;�R�x�oU,���VP�Qs�
�� U�yY�+�|����ω��X�g�g� G�u��'�8\@0�|Ԅ�������-�Jmh�z���]�u:�T�(r=,T�� ���}g߶�(��~�8y`�(��ͽ������E�ܸBv@�g����T��Y?+~Z��
�mvх2��Rwt�2��0�@��K�E��%$�F|����XeV��%���+6�ɯ���j �NY�>�����D��3�oB֬��L����6���많��x��y�O��Kպ ���� �O��'i��z�Z��2��HG�(g��Q�݊s MF%��㨵��v��0��/�ZP�P�Ӻ��<��'qP��LoK���3�啩mT�εw8�{!(d�Oq?`�c�f��k��۶��GQY����a#�鈊�,�����t�Ӷ��Sd���}���PZ�%��t��z����7\�.{��R��?����ę&�ۃB���-��e��x���=.ۢ+�kk��B�G_�YӳXXlxVHYEB    1525     840�L���0#8�cn�񽧅 '/[��6+/9ޔz@Ɯ��>�i?
�Ԙ�d�p��wi�>Z�ٽ�HD�+`����@d�+!������ ��S��

�C���+o��Ⱊ�R���8%?Sٮa2x�-i��Y�p���T�������U��|�/+H~�+��ރt�G=Q���SQXz?/�~\�v̯�i�λ��v�w�Y� \+��G����]|gm�W��X��7�LS�e��ߖx��&ܨo-�,-�e��[�?%Q�P�F `z��in��F�
�=�h('�&ۣ�D�~��.-����mX��jƸ�g��Rԉ�K,�4f%ż�w� �����_#y
��_e`��]�-GmR�<�i2�uS�>�.���m��)8�*2fh�rPA�!���t�z<�d�j9�/�X��m�֥Mzr	�)Z� w%�n����r�2+
��_�l�ޚ���=��I����Nnԟ�����f%��ݦ9�/�_1�Y�v�E���.
�z]t皪\��u����|�*J� l�&�?��y��Koq��|�hx2Y�<�V�[�˴E��Qa���a,{�`g�)�k'0�#���bf���觎�w�?�0�""�`:?���pg%��i��tH���B%�-=�6ƥQp�=% �I�re>�,�dأfWQO������B�
O��>�0���#�D�g��5F�O�Ŵ��Ϸ�9�#ynz �����K&��
�%S�ҹ^08�\1����.AxY ^x/��gȺ|�,餱�j��W��s�	@��d�w/��7�M��h��A��D��D��`�Vɹd�!еR��:�W?'3�4�^�ޕ�7�5y�R'���1�=m4iy�ׁ
4��v3I�����vB��c?yQ�?lF�����m���o�R�8^�5Á�?�+u�Bzn��ղ���d�)��ۖ�s<Y5��kOCE��"��o�e5"" ���~�P����1�z�f:�0-ke� `l=))sNE� ��%.�'9E���d�<?�t�M��?�4����܆Ss�SxYKx����;�2�C"��/��a��k(	�Z�i`����Mί�@���|&&\4е ��{�^Γ�:@
a(���+�g���4�$.�'>�cb�xv�I䬑� ��U1��Cm#O`k��Ӎ�ѐ�ZK�O���-���K=��b�RK�u�һo�YA7&'�6�.�Zx��A�^��_�Ԗ�VA��F�V#�2��I�=��i�nÔV�Y�@��O��������ږn�������Z�����|70+�\�W�3�h��D%�(��aqH�3,�hB}�Οߘe/�1P(b^�0K�f}a��h�uл'A���tP���KDJ�4 �'�r�*r�:��)
�D�̙�hz[s�=�#���h^QdvCl�_�4r�����H-����O�ڝ�akD�Ŝ<_�ʿ̈́��:����j3Y�]���V[�Sf���o��4ظ�u�f?�#���ҏ o��T�ο���l�7qb��æ���Y�B=m3�_�/��F��C����q��a^9��ϛi���j���z�Sa�ؼoU��O�&K�e�+z�ƴ�8�Q#?���EwG"�9��%˚Z��t�L	34�#������s������	CK��h�^�����6��aM��T?���Li����bjU#����E'�e��n(���nJW�ވ'(>s���'��k��Ryx��^����S�H� �vs]��ٱ�/�1�R@��0�d	
TL3օ.:�3�,�B�|���Pj����a~��|F�p�itC���l�P��<��jW��q�s��NŘ��	���Z$qs�G�&��Q�S�ԑ��bтy�%\=@��:cج��02(~��@lw�8� �;��U#�fI}���%�w�����\ώeL�<�����#�?]y��;�*�_����\���e�X���v���n�#|���8d�4��e�v���N�JS�	�t���ǖ�:5�>6�7�!%C��x����ïs|�`�l��WA9�;pz:\�x���˝8|�����t�����ev<����o