XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i�M���j%APx�E�?��F�_�Ӎ1=bZ	��1L�썊��5aW�g�_��4�^&J��Qh��J)�zFQU�,�[W��0�O��RC�eZ2�����ؼK������>��}b�nj�lc=ĕ5���u�ϳ !w&r���!�˲I�6��A��3�	�I�0�Dj�(���H�;�pԄ=��Y�G;v�^�v_���7&odTu�H@pdB�%�?���@��	>��[R�a�溚�#����V���DCX�'eZ�_�%",U��I�W��v-�KAx��(v�%P�`W$�fø5�ƾ��-S�]����W[Ѕ�)c��ut�����Z׾�n�?�]P����*Ϸ�<�qng�4��������ea������@!�:0��2��~���Ԁ�H[S�::+K�+�|��g�n�N�����-�dz�nixݿ&�,��3$�l���f��*�X��!�i�^��0�@'��y��(]e�FWV�u;������_��G���J�S��04��C{ �V�ƔR�?���P�ȷ�`f�O���H��К?�Ҁ��{�J��f�u"GF>�]J���u�\=}�N1y|�íQ�H�T�U=��R��ˆ�7�vؕ����W�M6�2K� �@'N��i��(�1���Z�:>pX	Ujb��yG)�9�
��Ub�n��i5�mᮕ�3��HI��8F�J1�}��wWb�UHa`M`i���};�Wu��X̥^ԭ�ϒ~�)�_�XlxVHYEB    7021    1e70"LW���y��X[N
��B#��ؐ'=���.���flg g�3'�0
Ͱ+(�bME���H>7^F-m� J��g����X��A�[+x"e��f7�ʗ�Rю�V��r8���� y�xm�/��V��:*4����g>H�a�B�3�dy�	�jJ�J����1�&��]������r����.�KC��[<��h%P�nm�j���=zF�`��g �8eV�|�@Dͨw������c,}דn�,��,%d����D�~���$���q1Hcr��:R~�y��(u֢8�3�;�'��쉵@w>HQ/��ZY�IuhT$&�-�Aܤ���\}!������XZ/,��
�wM�Ɲ�Ǐ��[�R�ωRj�^��<�.�����ą6�v��F/xv9��V\��;�A�"���gj�W��e�n�9�h�s%c��L&�Y�|?��/�Y|5�[b�Vy��-Cp6
�7ExLkx}�"K�ݧb��zP� $
�ƪ��ZU���EV���_w��f|h�j_UB��Xͪ��R��'&�-��>Q��!���u\���DR��u,�.��x�������ޣ��57B��!J6Km���+���aA�9u}UL#��|Q���j@�ٷ״����'�����(U4"��z�t;��r���N�m���B�M���:A�C{����	�f)<dc��p��i,@�4B���J J�5���������I	�
�8�wc�]8��3��Y2'dv��Z��L���"��pt�&��������F~�vQ���d���)�r��ٽ#n*��
��h+�>��؅pGh�m����l�A��*��\�F5O��[�/nԣ����!�Y���iY�@B�T�D�gVܬ�Cڥy�d/��$ ����9�2LL��V"zڣ�'u��02�hz񎆮w��\�؇�P#��;;]r42z��5X�d�.��"�������`�!�A��Y��i��?��m��$?�Kc{H����x`<��Ӽ�0r����*+)?�Y�.C�o�Ly�à(J\~|1#��kpN)_*?:�:{|��L`�J�9�%\�g��Ck	��7��YH2�F{n:M�>�uU��R�"����k�`���;���,:��ג�tQ@|�P	�jy7
��,r��JV�*ɧ]��@ɢ��\�� �VW5�DJ��f��oiO��ּ�XB�3�g������T|dsd|�܌��8�8����7���>�#���$��:4�CA�X����K���`�3g>���e�G�F�n��&�b��y������m�נ)�_�r�M~�0�"g�P5TJ�ż����?�ܒ?�#�yW� 6��=}���8�J��l�o."�e>�`"�d�\��MdSFϵ��1���ڨќ�@Ws)�~
�Gf��A>�����0���Ů�1X�3H>lE\����h�O�Km�$QH���#�*�c,������O��?e #�L';��y����8Z�ڛ��_#�w�	i�I����|I�T�8�����h���ZL�M��}�r���\m
���R�����ߪ�r>�O��\EY�e�Bkж���{��ɡ�n����a�@����D ���+qDu7�B�1\Z�T�����أ����Q�o�/h���c�ֽ#�c?b*vmLs�JV\\�nH�K!�9�2�?~�sq��v&��Kĺ��	V!��j׎5��7�`�Є<����F��\`��G;*�Q�X�k&L���"� ~-�ʨ�ݖx�=S��j��e� ��Gn�g���<vs�1�a�C��.��GK�C�t��,���;.��*TOh��VϨ�ֲ�<sX�_x�|���ݫ�^B]V�����y�Z"Yjg\l��ơ�p�5;���4�$����p}��6"v���a��K.
�s��_�8���/F6��}�
w	=x��n�v�#&��&jh51%֝��P�B�����]��,���bt?�8}=���,��?)L��E0��� j���W*����~�E�D��őJf�̺�9u��i�,c�3��Ɏ_V���7�݃-�yR�}�o�Z�P�O�2"��#HeRv��~�+��*��E��ZZ'�I�E�.����BR�C�I�FSKm�P��-Y!�8��O��>�x���0��X��Kl�hJ�����Α�n_�Apku�`����ɓ�'��	luTt��� ��e+]�ݡ�Bn	E.0l�ݧ�����ݰpo�GH����R��hs=h�đ����T����٧m�G���M�'9飮}���m�#M�������9*����D��}�/7,:Ű���`�����b���$�6��|MMv��dcrM ���'���[.�k�1�Z�w�De���V'#W&3:2N0�.��'�b@��WDI){^�
����}CߙB�����f�h���.H�a�o��v��%��E�ݐ�lP^�^|%�<7~��o̙�6Wh��d{���	��f��&0��#��>�'�>���8z�����7Nb��4c��o�N��1���$�m6��+:sm�u�$��/`��u�u7T�����)$?�ɤX�,�R�qY�	/���?��5���:���'dv�E_���h���ؕ�9��=�M}��sH;�áާ�OP'-n�M��og�p6�V9��J��4���ae��ɃL�޶SU�m�Hʛq���G`�)��&����-}�̥�9���@L��`�V.`J_,+�aA��*�C�+�Z�g_сN����c(6�ܮ�=��8�|M��P��$D�g+�~�
F6M���Op��w����н���\�J�`�-������7ǯBb�1���"hܶ�20�=_^s�T�����Q�T�5��ч@��Î7�l�� �"�?8$��t���۩�l"�t��R$�a�i��L�<�,��P��#�\�9�&��}�72˸�yJԙ���hˈ�m���My(GF���֨Y�6�<�����^����I�OF�2�d(��v]�z�����dN2	���|�N�DC,�%�JP��!���f۾������`��W��T]�	��x�Q�bbW4��Bq`ͭ�`��D�����|�y��@;u0�Q���"�	��
��'�1�J�`X|�O�I,p(�UlЭV�e���\)�(�O��{�Y�[-�X�eK�n�~�����b�h��"�+v��X�yy�IdBm��it]l��%�i@��Yuy�&��l�m��YՎ0�f��R���H��z� {kr.ŭ;�ɡv@�D!��&�FaM}�Il�idvY�~/��ٛ�P���t,�Ä�]RI�-(C��<5�'��L�EVY\R6<�2V�2.��.��/���?"����oc�#9$�� ��p�%m�I$�����W@j?����6X��ȸ��ُPO�pЗC	t�V��8Y����.���ab�ꤪ�L���H�X/�:��/��b�)� 1��~�pm�),"wl�L���Y�����OPє�োx�i�����3Y�A@���K.�r�r��`z�OQ����P�K�����u�<c�@&�ԏ���l��/h,-Q�^��a�t��u�~n^ֺC����kS1�;�i��/�2�.[N'�0�6��s(_�`g(���%�h���ȟ)~�7�f��WR�'8]O��yYJ���&��H��!F�9[��P��)nPȹAA�ðc��$NK'?��l���(��Z���Rc(_�]���L*
%�7�-=���r����l���  sJ�~����x1�=?�M��i�w"*Ԅ�2�����������q�2�o�q-�@�i��1�3��X����C������l�9�̂uE^�Kyk�v�iE��a�0~2X9�c��I�k-F쓮��|��>��4T�t�U�w�&��%A?.*4
���u*��G1J^���",_w����#:���L8KlK-���Vg��	���;��v@|I	��P��t�������g�����*o��+�B;�����r�8�I�X8[��L`�2�: M��S�=�_�:vJ�S_��/B��᪝#�z)� �M��5�~��	���� �3�z�$�7�a��Ntq|-����_s
���l�QXo�9�r�9�BQv3���I����$�� �dcvN>r����|A�T���[�8v$Ubϱ*��y�S������G�G�p9�\��ԉ��
�T������K���c�ә�����o�r9��M�Ͻ^<o3���w����'��MB���5�l~z����7�	"��f�7���ۑ��6x# ���/@u�>pi06˩�'�I�P]y�Lvu��)�J� 2�	��/7|�|7�`8�C������*r_��=B~�~��i�E݀�H?�!����U�cK�.�=t>w�D�������ڨuY=��*"�Ii���4����¤�Q���*����V��.�\+<Bqn�q�'͘I�"����2�8�cʃ��DS�ö]�f�[����E�|��<�'s9)C/��|�R��̅�>jX(�锻8�(�_�Zba�0���ё;Vk�p��Bm]���Z��ڌx���-@A�`�נ}����?N�n��ֈ�L�QR��\T5���}i:�Q���'��	�ƪ[/�V����x)����L���\���Y;d�
�m)��Wـ`�[�����Y}׏��zO -�,g�ֶ-<����]�F(! ����#Q�}� ʜT �ms*<L?&X��ը]"���&�d>�&47c7��:��Ӆe�ɉs�4��+�RQ���sfx��`H�Ȁ����d���.�����K�T�e���(G6H��g0��`��g��QJ�;1>-J׼���dM�(�͖��P!P�SW������7��G	K��	U����5.�`����UzJH�z{�ǵ�9wS;}4S�A��^�w��{�RO�����,��형��j{NI�����|�Փ�d�;p� �b]vp3��T� ��)K����P��AB�t%��>^,[�O $���(z_����K�\�9Χ�P�:���_'���d�]���[�m�2�"r���B�VY	�B*~xP���[�Ժ��j�l
m���臠�R�)�=�Dc)YF��;���JS%f��;��B*���T���;��&'8����~$u�	V������b9)�1.�F�,y�`�̊5�(Ǝ����IZdtM���Dۑ��n?hw��=`�k�Q�2�rߦ`'��e��f!��������Y̱��OX;��x"@؉�'�4ͺ�OxiVS���S��O�Ϩ��޷��hWL��x�7b��"L���@7���C����4��]�[O��5�cKO�K�(��čv�g���7�cY��Xy�F���-N'�as��q-�<�'"�XgAk�tIp3gZ����}$-�MnZ�?��܍��A@�SPZ �=;�āoiH�EL��wEFD��|,b(��x�Z����0D�LW������FK椦~#����ezh1'i����0R�*�W�GS�J�Mc�PzgX��5���P糛���:�����M<���l�2�t��̗���R<�a�G����+Aޔ�ES�хY��rj�b�L)s�7Qr�.���9���� @2P��V�ݗ\���_v���}��1�7�'�~�~�s6Vᯈ�p�WU�<s�1��1����l� <U�B�%WI�al�#T�;+h,�&l�8K��a'�z���x���I�8���ѥ�R��s���S�|N�ԣ�K8H��l,�\8�횼/�\O��7��T͈�V��^�4�x�u����֎����>��G�R�k�o|�M� �A��mb��ѓT�U[��y�����7I����ƪ���l��A��R��<p�5�v�I�m+�T	�g�>/�M��ׇ4�Ԙ�����������!�Ԃ9���ӕ�?�W��)鴱5��v+��$QH�ϊ���2#O���i @D�)
�'3�p�j��'��ND�	��_��ѻs��Y ��*�h�~6�|��-�%V��oR�)�dQ����+y��R�ll�5ૣ�oYe�s#b�3�~\)�h9��7+B�] /�a��d�q�i5��8�!%j�nI�MVR_~gZ�n�Պ�a��^:�^��bQ&/����-����a�Z��T����9$C���g*i��B��~��$.���oZ U��C�"���/�k9���//(�eF^�=Ig?�^*Vu@��l0[��Ҡ'�{a�ʸ����
W�.p�:W��=��QR4j�#^Y`�AK2��þ�¨~�lᵰ,���U����U܆D���"w\~Uv(�͛k�G�oҏ%��R��"l�z����g��c�,O���70���h^�*�X1��0=����Ɓk2"���y-���+�!���NX�\ ��t��(J]Ox��1@�K���.�����soȒ���wE F<�7��{k��ݤ��-��y�V�&7�<q�:�-�N��:�(d\ {��K�e9[=�?�;�MM��L�z�S;v�~� �i�9m�&7�
I h���3�65}��!��-l�͂7��k��=8�L܌z^�Hu��D�Z�!-��;\M=���\���������?Sʲ�ņ�����׫q�K�R��e=ҡ��
��a���܉ֿ���+��Я�h��O>���G��z���{��x����0�0�9�Ȱ{jMG�)W}O�gG���Y�+۴��YY��b�\�,b�I���ĪߏI1'�YG�E���1Q���̄HN���Z�|-i��^ǵX���k;T�����zX���i� =:�|)y�Cɼ����nh,q�|�r3��[?��H�o��m%�6���b̚������j(n��c'XfyJ��[�Y�v�~bPe�i5#*pȡ%���׮�œMԤƬ�h�}|��(=Sl%Q�6���81�V�� b�8O6of�,.GKvn��+q�g^�������3|V�t���d� E��"�Z�*[]�y�Ph��M������o d~�r�e�[��8b�0�~�C��q�m��Ţ��|��V�'��[��跻y@1���l�c8�sf��]��}U4����٭�"tl�"���Z��j����q�9�u���b�#��a������\��S�2�b�
+��$]�$�1,B����{f�v��mS�������)n�7��H̤�g�2d{����t��IAwS��O�*��O.�g�wN_Y��)w.�^ ��}�|w�X:d�Z�~�� ��ʆ����J0�Y u:k�^��Ӽ�DԦ\O���"�<((��>�l�&6!iJ��6�n�F��u��f��:�-^��M+�jٌ���y?H^�����nY��\}�ŷ,Oڏe@e2<r@?�w�O���d�.ȯ�H�\Z #g��|�c��(]�]|�$�*��,��>'B���2@�#{8o�9l����Jhc�c;�����ݲ��:���Vj�f�SC�ۣ�1M�J �S���&�B��)r+fM\BB��MLoӡ�����/��g�C�d����p.�|�¦�Z2}��,�Ժ��w
�O��"����t=rm�e:���;ϻ�����?�#�lW�6/��&��=���<~�@��,k=>�;�:�\fIs