XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ې��
|����%�̈�%Uc�^������륮�9u�<߸IS�G�H6�@�:�����ۉFH������8f�+�$2Ԕ	�u*#�g	n�,A9O'����f�~:�V�M�>w�.�/f1e@m	݇G#�.�r�f�C�8 u��@a�����)Є�d(�B,��a�CM��EH����O/�1���R:>KZ�.?���Q*��Z"�����g���
3�6E�	R���~7��֩��"^��S�A~'M��@Vݞ�C}�������XZB�M�K�R�L˙���]��c�Uڲ�S)���rݩ_�y�a���B�j� �bX
��SWKU+�l��2ؗ��;	n�+~-E�e��u�3� �'����>�Q=��%/?JԾ�}?1GO<<*�(ǛM��0���k7+e�ֻV����'���1I��/�N['�`
���?R�-�����6�ԙQd�	����C3n���b�GRYa�O�~�²|]qz�(w6�Q-�jޮ�3��铹6�'??�
�ϗMGk�+���K9��9�x�E�P�<�Y]�o��o��jy������s]��S���g�l����9�"7�g��=�y?Au�v'���o��FD�b���8p���7�a$��^�ߜ�xԔ�j��`���]@�-�d2>o�����"��72W�N���h�|��I����d�d*~�D"�<jx	\^����a���hBPuV�l��-gy�����?����B�� ���#L2�o�Ò�K�����XlxVHYEB    2d8a     b90~�ԙ�@D�{y��!��N�PyU#5s)�~�=�8MqA�{�!#ʭ'�9�+[�i�9���f��k��Y:m�*�Π�����f`l�pBq27�B�(��Y�A���q��%+d_*�H���z�LGG$���n<��:�}��OE��DKI�=�������[��.��!N�P���s3-��A]1�Č��QI�U�aŷKe���5u�(k�_�)~���4��i�R�"�;0K���dT�u$^)$�����5���hO�����q�&m3aoM��~`?Ǯ����G]p����3$�����Yn���P��e��l:|d�~�7np��g�|�e�4�M8���rn?��{N�������AY^d�!��a([�����
�#v���5Ȝ_��̯T~�@[:2M��d�jA��c�z=��T*����M�vaόw).B�����I��z`!����%YSi���;F��,���e�������<v2���P�B�eӸM������f����{\��jI��� �@���OgeQ�'S��O�M(��ï#�M��+[e^rc�9���y���k2盦���d%��q�ǁ��.2�r'z���Fՙ`1K07຅5������*Y���q�C�]ŞL�/|	�CB�g;�=3B|�O���گ.8��5t���q��T�I�gl.����1�T*���TQ���D#�n_�V��q�E?傪�뉥�|D5vl�TxX�yE}#404{�W�ie�(��/2���@J㵕�Q"�F���A 2�_8��3�� q���mH�XƦ�AsП�P�+��nu|����6���ؒ��ad�s�X0i ��e[R�4#�OET�~Q
V�
����4��J���'�7W�¸�H�^qSBO���گ���O�(�q�ΌԼ�1��[�Z]l�!�eY\��M4
�:�����"TV!H,���ټ-gd�_/�T1��=N�+MH�&��I���5�.�l�����}�V�ů�pͼ�]������݂�FF�u'�{��� �����@8��(Y�'.6��`��b�{k�{\W8B_�
�0���ΔF�β�)��c��H��83+uZ�u1��{S��?�I*V�ǥ��z1�Wj�v�W�@�Y�T�J��h)]��{�'X��s��R�)tTku�N��P1�c^��)�(݉H�A� ���;�G۸�]{x�����ռ�o��C˥%§�8=��WB�%��ȫ��|6�o0Q������E�C��D t��s*e�S��=s�s3��B)Oƚ�hŁҚqeK�G�A�iu&��6UJ-�W�)F��`�̾���Z�����p?������U���i�{]��b�����kD���&o�3l"��۟v��{l9��#�
$�^{<~Ŗ#Tfk*0��&1A��p�&�/��K=�_�����+�м��#��:�D}�GZe��Z��><�-ƪ�H��]�R�;�9�i��T""��O��AՎ)ҭ�'���$�ڶT�~IZ{TB�3b}/#r>0
y�ąU;>V�L�8�E�گ| ��b�`^f��-���j(/��#~h>���e���&|a	�k���6�
۽R��h�!��<c�2#�M�5]yU���w��`�t#��zT
����j�IZ_������a�E���!�:����/4+jB?�Y]���d�������Sk\���}YKX17~��P�PՖߙ��'pk��ʖ<2T+4��f)����d�h�os���,
��������=���P�+��[�r���l����Cɮ�u��[��s{����wx�@��xw��#�^'ӷ���VȜ�g�@ʁ���������(�.�%w�4�c�&�������Ь�G�o��"��b4L�bQW����_`0�hƀ��S�'+h}_O��Z�[����{�˳Z������EN�m�run�N45XD���A�+ӫ��������,�!��8��Q���D`�����g��7;� ��Q�p���&��yW����P~8��ɟ��B�AwwS���V@@��/�v���<D1НM�9���FRw�7e�2���~��r*����\	��S�ŏ�8?�d�c��P3�g�����g�`5!@�sw!]Id�/.ƅ��6����]CA�gN�N=�)֨qm�
��B���T�,�-Xwa:ܸMI�lQn!�m;	���{ՆI�*���I�lcΉ`�����⬸V�G�艀OB�x� !�ډt��W��ښ�EHJ:���1cr�Ԣ΋�_�j��Utܽ�zZ��Q>嫙�����y�C{",�Cn'�O��
KŐ�����ͭfR�{u��/,�O�(�@ߑb2=��� %2��F�	�_5�	�TU���3���)��c�������OO�����&2���5u�Cx��>�A�/�:/^#_q��FN�j���pj���v��x��tV�@���a�jt���?H���8��9[�+D�Ju@�h�2��ߗ&�
��v�*��΃J@t3z�ฌ�����'�F���CvhҔh<�X5����`D"_�so���s�+�f?�w0_͓t�)oU`:M���(,��hrU z���ă��K7ˣ_��N#՞p�������r�R����D|nc��7 ąR�N��"O��0�#,��O|l��`}9��LC.4@~�~��h���n]o;�Q-^���������q��(Q���9�4(�r������s���1ދ��&F#z<��w�N���;�7Wk�\�O��o�ET�P�C�u�-E=Kp��4��tA,Mo����z��P�]4�hc�rS_o��p���q�7a��>������ ����Zӻ�#��+��eE ���A����j�<��B0[�i�ȑk�О��Z�8�B�I���tS��a�;��b:�s�Q��