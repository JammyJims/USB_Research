XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������W������j!=򵸊��|��Q�^�9��9]��%���k�|�e��Ng��]<4����{���e��������?I��Iff�,�C<@ ;���b�M��6�ѫ�
̖^+9܄���J� �D�hc"w�M�/P�R代ս0�Ozd6��E8M��e�~"�+�l&4`��ކz�Mz'Y<9q�P��rQ�K�S��hf�b�d�I���]�(��%��q���t��� 9�Sb�ǬY�_&��ޫ�͇�#l��@��E=��?Ȑ�Z]��u��=ޑ�T� �Y��9�Dbx�a�"b�����<���	C׋+>��Լ��>�q��:Ջm�}�oS�����a��;�Kd��`W�$bT��	w��i+�m�#����`ݼޚ'�wf���][�t�������l�T�-oAuv���R�=1��r�\_�04X�W_^Q�D�'QP���D�晷�(�ᶁ?�����a�(Z'��4X�I�k����J���<O�B����#���zC�{�b��y:�皉,\�-i����zsA/���ccg��˺�w"R��T��@�~ȜON������-�x�\�i���J.��~�<���7�]����'h).��b��ꄍl�p�t�o�ϫ��ˎG��+��Ыьl�<hǴ� ��Tv޲���a�j���iߜ�*���b�[��g�]c�+Q���
&�|��=Ipҹp�l�E���4�XlxVHYEB    5103    1760ą��
�w��c�����귿��rp���}u$�
����*1EJ�l,�=.��Q���Я8< V��`�Z�����?S7���xp0���˲G�\W�:<�\T�x��cM���:d��}ߺ_�ܜ���"E�-�0�h�JL���瞨�a�Ƣ��ܮL+c��H���/��l���[��6�$�\ݶ0r@"�E������������������!]����D��K�O������V�$9���!9I��󚉽�Z�a���8U�I��#f�3�kB��_�M8H�N���R9i��d����%߱;/K@@:�]v�ẝy����?E,�/�� �Z8]����@�fչ���7����[�������*�ЦO�{�j�h�!�������j��6f�̺��uf�Xx��т��#�f()C��,��G�UW�2���`�G�z���:������)K<��LXr���EΠÔi!�Z4�l����6�� >��4�ɹn	���Z��7�n�+a�.�m�A�@(GC'�&���]�4h�YDt'���8�$�v�����x��k����L@��p�8`�DL8�Fr, Ҭ�98��
"dlr+"�8!'�W��� ��#��cb�l����ܑ�� ?�W/�ئ
�\,v��cp���C� Qb@���1�Ε���z���T��Y�g���x��+���y���]�F.$�|d��d-ʦ����ШЏ���NPB��v`2�����PE��3���B)�W��K|(,
��#k/�����d�*��l�� kTxz���9r'�I͑�X�a7*�F0	��5�E�������C��`��Q����O��$W]���Q�s?E��^Kv�q�^�-�C`B$�]�)��N�qN?���Ŵ|�ħ�����rY׃�ы�q\�1���쩔���N'8|�r�b�����%K��7�:
Hr��Ǜ.�T'�S���V����)�Kӝ=�D�M�i���b��Iz��pN
��k��d3 �Mn�U)�y~�t�p|#%pn����tPp-ܺ-DƮ�a�;Q��9�I@ׄр�����Y�Hk_p��Ć����/p�c���щ�nVSpP�����A�8[
7�ҭ����]8���u��VN%}^&)K�O;o��f�ϋI�@�"u�m��)�p�ݞ9���NV3��봺� �@4D+佶�Q>37�b?����m
"����	��� ���k<<L"&�
1@ܩ:	**�	��Q��HB0ڶjT���c�_�~_��D�����*8+�O��}u�T ��_�[!�P��u�X��"vh_��%/���#���qر�A�[&��J�
��"�P���B�C���50g�����{4�K+��ػ����G0�gI�3ce�u�t�vq�v@ؖ(�Ք�B7�<k}���s����=��[�}d�T�*ϗᘟ��R�SB�����X�?�s>��e�3�=�j����]s�5�xL���y�N��94��V�����Z�ɮ�=�QTˌ�M��u��1�C>
�H2,t�WYu�/f�숴���?���������$���Xi/ϝ>>@�<�4n+�徭ĒKJ�s~\���Z���
��۫�g"nv-e�G喡C&v��y�菀�V�! ��t>&��|`pX��"Tsh���o	������-��)�H�{3�d���$��cX����Y��Λ�CT�zYȮ7P5�$9�v�NB�0�Rf�Fu(IY��H#��\���i���$�ʄ��B�r[�~5/�G�g-+2�VJ�`�3� �S�'ȃ,����>r�A?OS�N�Q�.�� ���*��kI�B���w��i]Á���|0�c?"�h$�xj@�f��A�q0px��]T24�C}�κJu"�j�F
q�mJ�0}(�<G9�w�"�O��;�|�HPx)h��]Z�Cx>7�c��h�HLv�������φ�{���[4}�2�;�f�-�,Ki"�1�_�%���<7��=����܆tyW(����?���`�X���s��^���h�{�^y{˃-i5y�� _E�{���N�	Uق��h�^�r7���k�R&�H�?��Q�L1v�?nj��J��g���h.��:��2G�;)�� Zɑ?��Xy�x9��Z�~HXɸ8��@�q�X�8����.+��r��k<rn��s��a]i'��j����eJ�w�
�d�h[(�@�W�Û����i�a�C�*������{�s=P�w�	�r1�jtt�P�NU�F0f[��\A���IM�S� ��w���كKa�wF��vK���JS�AEm�a`�8�.nbe��g��{�3x�2�&W��� c�3�8�n�Wm���%�?�م�z�Rl2��؀�g4�5jw���v^6���ì�	M�^�0��uPF$�}K&�Y��W�M�B�EY��������hԁ��������2ET>bH�%m����݅Q:���T��� g�s������G�sarR�hۀ ��%ڎ6�y�������F�����`�v���~\�~(���*�F��OC漲��@+��� =��><���h���dw��[}�ـw�s�i��w5]V�)0��ئ�\GFВ�}mzFQ鴳�'�Z��Y�B�r���uZ�Q5Ã���^���+h{"./�:h��j��~���{�0������^e��ST����쵰�� �Y���>�@��B���jɖہ'ަ<>��K�i|-������h�VY��<ǟბO��/2��o3�p��zh����-#E(]cXX��+�A����]����Q$�z"<�eEPr>�R�?�.J�	�MJ��^�T!z���aĊ��Zh%:h�G��-C���S������|��S�P�n���mhY�y(o1��=��$�ȃ-��3_�(��N��
8�7�8P�p�0����
�����N	A�Ck�ň'�<�6�]�$<��>X!�:�:<p�����?�N1#��y#��$&��˕��r�Yar����P�˺l�l�4_���-�+��侱��!���tj��:^_d`j����L�e��:f����7r��� & ه��h.=�g�˱��V�� Y�c����bT!�<;��WF��������L`�$�'�:ıp�'��L��~`�_�S�I6n���ŘGS͕�y��w�_����E�@w>�~��� }���y���Z�6]7����S��L�NUa���Q,%�S���#ؔV�f�'�
S�P ���{��W_RT�3hE?���������
�_���.�0h-�5����L��܎ � �����ځޟ�y�b�HD/�O��N�[Wx�j'����9bǥ����)�#��D�]����.y_2����1S'����?0l@"�7���<�ݭ.7qm��=j;bO_�(U�*�Y���|�}c��],t��\�j1�U�Z�<eŪ���	4�B���C��������7~$b�x[MM;(����E�c���bwK���@m�n[@����/��A�!�ù���!�Y�W�d]���:��󃮑�棌:G�V �
�J�ƌ���~UJ����[|�36C��Ms���2?y[��8��5��$o@���cp�-^���ǡy����rH|y`���5����y���Uw1b7 qE#�;!�Gߍ؆�K,/��HJD?�%���6�. fP�h1��rY����i��=��-��=w��^_qM�#�s Q�L� ��	���x��!� �`�h��jg������d̡�?�����D9������bb�<��4�a:��\[Z�kj-�� �Ԏ�n������\��e���W���=;	(R'�$y`.��G���zܜIN��*V�L�W�8^���	�Tq3���
W��E��²�Q��>��.\S���7,�#����#<�.�&�W����wk�d/����=��L��{�ٞ-�ʭ��U��u9����<(�K���O�D	x�C��x ��$ﵨ4��e��3�/Mu�򶎡��4�'�{�?BL�_��>��?�o^(  �v0�����2��5-��J�Ԗ"����` \�H��M�ㅭYknoY���m��@��x�y�c�+n�c���,ҕ������CEe}g�w1}�� ��L�Ɩ@��}D\���zr�����������eg����J�7����Q��9�a���.���b˽v��W�^��lo �zn�}�d>��!I%n�d�9u�"���5�*YfUIک��T�HB0@|: =@�=w���fc��������k�٨{�~s���ǥ-6j���`�'���W/�|r��r������Z�Ko �s�"ڍ���>�/Q����(��	��zP3ȧdu�q��` �S_��P�w����+|sm�~�w/��&�O#�'袸��VFm\
g!#�KK����D�6���U?\�{����L6������ V�я�m���I��{]�x�m���d�^���9A#���Q�l`C��足)4� :Pw��B��XǱ��M�l+���$�J}˞b0��)��H���G�[�� 
=���\C�z�8 �k[o�z1�In#�O�FA���bS�삑�2V�$�6T7�(i��Vr�w�k`��]�N��c((���̪Ǚ�~�}u��Lc��
R��^P�}�2���̑�߂���������NQNXxs��󿈇_�D���D��!&��"�����^�]���"c�;Yx�A�a��I$�����rQ`�װ��k�h1w�2�¹#z,��y�I�0��a�V$�O�ފc/����=�C�%c��,	9��f7�VXz������/�a{�CA���.C� }�"���0�X��!a��N4
�b� p�	�`���|7ϱ}�뿀h��P�3f�,
!��S�\�Ѭ8(o���f��ї{��YL�I�x��nGV3z�iL�����S�&>i��b)į�MAv�g���D��>nd
>t���q�_�F$��44W]Z,<Lm5wx�4j�䓣�j� �e��A3I�.\,�F�S��>$��Px� :����6v�աkt�ș��T�ķ�*/}CX�!�/�X�H�/�e�n��{�P�]� �ѝ{�eS�71.�OZ�n���gN|-�-osj�W�hhȥ�m�����p�dEA�	�2YA���\g6PҾC�����������xq*k	��5��aj�02A�.<Ч�?�J6�~��C7Z��sl}�Xj���XF	���>�x%�Z8�tP���'\K���_>4�LR�J�`j������BO��W�*�=�,&��o��#�p+R���Z����	F�!k8;���W��ftxJN�4m����e�v�ؤԎLlz����t��}��DH�)q)J]n��![�WA�#�^C��S-�qDa;T�xV��H�4�'���e[�u	��=S�Ub�>|ɖ��s�D�� ��Հ%��\IZ������A�Ssmן��������#�%�^Rr_�\[���m��s�]��_�B��sM��g�\U12czM��b͕ $::��N?j��&b�M�b��ࡖ�vs#c�U	O~��+�'G�@4.M������R�B2�
�t�ņ4�&�s1@wsJ�;,�;��:p�?�v��֍|���(*/����D�Ӹ�7&�w��\���M�(��DxI�S�F3���y,�����y�|����?�M��d7�Z�`+���t�>�B�i�����=\W�K���&��(���_$_��l=�0�K`U��]�f�������;"#d�kX�������a)B�XH�WBԈ����(�1�ƪy�����^���3)gi