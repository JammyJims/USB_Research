XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\��-�	5|����㚔��ݭ"gZ߬"�6�L�&��u�$H���/�3�MqQ����p�p���S�=�V4�YA&R�����er�I��p�?��j�!j��^^�%��X@t���3R`�:�jy$�1ܩ�!م"SV�@9A����8�u�f2|��q��b��55rJs8!0ӫ���e01>BQ��h˝�^�J9�j-V�=��5��y%���I�_�;-A�^ #�3\Lz��&���g�������b9�aJ�m�Ci�n2J$2%� � '3��
��>F��7�Y�w�*�`�����ć�S�����Ұ����rX�'� bQi��GhuWg��ƺ�֧Co �`�׫Q$A`�(X�QRD~ƞj�a�j��s^�7�Ǘ��s-���A�Ȟ1(���\���H��Afm��&t7���AP��T��3F����x]�����������q0j��w �j�[`)z��۩��xy��T�Oy�������!F��>���Kx7� "0�H�Yk�0��(����Ac�=9�q�S��3FND�!&ou������'�C�_���e��E0��O;e'��܇�,�Z��|ZK��?�+/'���̍f��nB?����S�/h0��24�%���;�v�[�cWO����KTRn$Z*���]�+�'T�S�[%f{�O`�2n)�J~�,����V�`<���}�_��;2G�/�z��i�����ZdʤNT:"�م����Ѹ{�ޛ$�tZΐ�C�XlxVHYEB    4797    1430^���I�ͺ��˛���ۚ�v��zHg��}}\��h�s1����F��p_��ԍ����0x_�qc(}�	�1濚�����^�K�7�Wf�H�$�#6��w��~�ٚ�Ǎv^E։���-y�ȴ���S6#U�Sg�3�%	�Qh�Xd!�a���p���ٱ1��2/�V
�I���u��;�zsU�֚P���N{�����WڄU�]J���˼^%����)���~a�jS��Z�n�@�$��u�A$���ԇNԁR0��&d�]֣�##���f���m����a���x����P�J�.{%�E7QVs{V}t-�Yv&������X�q:l��>��� ��^���vڞ��?;~tqS������mC��ý]��v����Eύ�#�;E���d��D�TU��׍��3?Z˞x�3�v��dc+s�Ҁ�UMf6�����X8-WPôj�c�?�'�W}�b��.&ky��9C�dW4�6��\�"A����C!��Dʇ|��&��'>U��݋�d���!��V}7Q��35�ء�3�2�X�>q4��(tLy������������ 1Z�,�O-�Å���W�����<Ҵ�tw����^�k�%s {�#*Ώ�l瀭�rD7�Gncs�1�=y �0 B;ϡw������me�fɾF���@h���l�VZDa�`L�>Zދ;_9��HY���`��ɛ�*����"�ŵP�yB*|a���0������+�;l�=��b�0W���o[�͍�n�.�@�x 3U�������%x6ĥL�˖�5N�͒�P<H�o3��^�T�10�As�<���HsQ�϶I7{�h�����yx�Gp(ec���e?xcC0Q��=�t�a��Z��(��
�Z�^!o��K�
nfMi��˗�l�Y--�S��Lp"�;���NNܦ��{��p��;�+�g��"�@����� ��|`B%5���Dב���Ug���Ǚ����B5T��B�R j"�	l����~ޘ[��-}�<�`U���G��ϕ�� �jwF,�,&gp��9�U��=���g�(�/<���8܄V�.���M���Ho6��	5)KWu��͹��v�e����{����U�&�aD�a�Υ,B*7 Bk���z'����aPH�fR����-K�5K0
ؘܻ�
���(������)�N����=#��.b��.s��μw�3#*�E=<wP�*���JaR����22r�-V���
yդ����{a"/��xp��w��s���߻����=��CXl������nhW��j�GL<��Kו�%X�,�Po�K�޾E';� �"D�ʌ�q�7R���[��������z'J��툫��R6�ؼ��̀�Q.��W�i��zI�� vO��"TS��ኴnxS����jI��W�u�GQ��I���,<�q���LɕM	3#���з�o�.�E'BB�F��������t�>������:WP|E����6��&����f�u,Z/���y��c:5�[ ����T����E�^����16'́� �A�윪�ѝiw��{�|eX)%�S�IE 
�K�������S�F@�J�J��ɢJLz�Y(·e��m�3��:���fs��N���]�q/^���a��=���t�·j�C[���O�n�H�Z늺��$���K�_��=�H�0�����	���ⴗ�1�c�ՃL\�<V�i�U�kQV�
p�#��P@�,��[�XGՑ�k��'�/k�aΓ���H�tflPdF�H�Q�d�0�(�f�X�	��q_W~�E�vp�]+^UgU�_^;J�s�E�F��ڋ#"�/�)��_1J �ɤC�/����3b؉F�R�e�t����8�iv�f�gW�L��Ol��t-gs-O&8`_%v����=pL䆐k��$Udi?ql� �%͝�V.��1*�;4\8�O�H���^��(�䴶�y�LA�L�=�'�������q�r�1�
��7�ar�@;^#u�J��Qٛ����\e�4�Z��\�y��r�|�w(�-��]��W�/0cZ���%\���~�e�xc�ӎ2�ɢ,�1,d���(���7�_�d��jw��&���0������]�]xZ.�|Z����@󺢋8q
�QCJ���`L�k;&��ۏV.�аeŖN��� �6��'F��Ia;3��_� �K���h�g�	��N`�ۀp$�\�V�|��6�2�١���'��4���3�<81m¥����~���b��N�P�� ����{C�#lY4���G�%��QYȥb���i�r�1���-��]����#��sD�Z��S1%e���J(#���M0�������@��?�`�p���>�Y<���7z6��f���#_<��+��x̮v��|�;[�0$B�Y����/-�:r\���W)l�c�r�#�����'6컷1� ^�]�i��g���q_U�8uD+�S���b#T�?4,X Bg.=b�O�i�J!��MN`@��y���:�@kwb����>��/�	9x�;�W:hm?L�/D�?n����S"r�P+�!���i���'�:k�l�X�FQ��\{3��|J����=}(.ĕ%����,A"����h'����KF!�N����(-��hkX�X&P���x�����o�	�䵪b�/�b�#����E�4>�uu���M0k 9�S���D92�E{LS��t�9���P�q:��v��#��^�!�*��$l[<���v�@���?@;��U*���eR=���Y�s�$1R��$;�v��L�P�>�4]p8�wQn�U�}��#-+ܕܟ<<mg-��?�S�E���;8k�)	x�����K37y��/����3r�]�lYpY.�\LN�nV��#�8�Ӟ�b�ྉ��q�{&i��w�0���>2�9��������h���W\��؆��v�G��X�z�]GP)�86�?����"��j������BA^�<H"ߴ-@rj=����	]�OPk��8�c��.C�*�M����R.-=�J1xQ�0�u�d��Tn�}������������u:�o9����2�3	z�װ�	3]�e�"�&�5w>x��{SIbE�N�GѵP^�����l$��ʫka��� 5Y������gH��E���d��(1�Û��M�q(vX�c#�L��4�.��)�g��@�j���V7�&�-���5�X����3YQ�ak������f!�Z����!Y�N5�W]� )O��kj�"��F���aa��8m�}��J��ń�!�%�V�[�eE�@�Fb�8�*���﫤To荒.�P�A4Z���b �^�Ѽ˛OT��\u�l�z�����h�B?�ۑ��tな��a�koh�M��!�=�g�?�P�-m|:(����C?��΋^<�%��5��>�#!ց����MLS���f��Y68R�'(�
�*ֆ�����v��?B��y����Sh�I%|�uT	(�?Y�a�D�����H�*����މǐԭ�qhߢZ�A�ɏm*�P8;��x��,�F��!jnH�݀4Qj�j���_��>2GHǷv����Yŵ|�_��]��e6�.���Z&
) �#{���n���W�H~��!���p��X����k�BY�sg�G����C9��d���n��-0?A�sӳk�;+��}`!�u��Y��[͸V�J���œ��S
X��7�C�%=H��p^����n�"Y+g}�R�"��9�Z���Ħ�Y��Ng�1������(gP�>�;�
N�^<�^�W�����:e˶-�O�������a��H�t��\3�-���c2��4���C��d�&5�_O��}�-~�j�kl�8�%��[\�d��9T���ژ�A�6��!�/Hm��4H���"4p#hX��A �}�"'�gvJ2��_Y���N
4����Զ�y�[dˡ�J���N�ê1į#p-RI�kOt`�6�����W �3�ɇf�`5a�"T�/�ʈMO�-`+jy,�����$��;TNL�[ߨ�3q�RĒ��Nq��'S�ZǘJm�����*�Ǥ ]u�ȝY�ߺ�x�����9�Rd�7�BxG+��V��fK=Z�z`I�T$��'�5�l�"NE.S����
��Zh�R�,D��4�1����G��س��6ԅ+_��;Nȏp���B�aδ�� �E[��(�f��3��u�S>��W"_����R�y��U� JИ��}����q�J�[|�r��T$)�oҧ�n�Z�&���b�B�wZ�2�=Js���-Q�v�`�E[�=�����%��$;N�����C�A8Z�w�\�~�ɩx1�}�z�4�k&j���!@kw�����`����%�=��+]����?��%6��S�V
�i��Ghap�h��[�	'���]tFNR'`f�Cs�L͞^h�T��l�r� ��2�rD��X����_�s�WNw����S�Z�N��zV�������Kr�s���ۢ��P�T��3m�}/T�չ�5�|���(G̯d7�o�F�3gb�������R
(�R��.e(7̤x�	���O6��>�&�B�C��w��>QZUc�vE�#Y�$ͻ���6�Y����W[��`
����1�	Ǜ��?�]ʏe�
�����+,X�*�v/{�[|�p��	C=� �L�� ���CK�e�הM���n�p����qp�$��a�m��tGK2�����Q4*T�N>R�m��4��K0ד`��vJcH�ѿ����2!Ӕ��mPHa=��!
a:>q0�ܗ�/S�����N@P2x�����l�dQ�K�k�kw����ȫ���)|ß)36�	�"�)!��B�&�&�L��p����A�%=��/�w	�������7l}^uھ���~�}��V���nkȩ;#�_ 6���G��(�\5]Fz(bY����7w1gŕ��*9�����9���W�:f��9�Og��ɵb麣�.M�D�S��,��������K$��e��	5Q9�-<k��~}��"��Fڙ ������1U�@`��4