XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=�f��]����l��aȷ��l��7[��
��|_�6	��^���=�6�}�HXEU(�3	敿���V<�T�dӍ�/*̯���|B�9��`�+h�p�7vd�B}�a��j���Ƌ���Q֥@Є@Ǩ�1���F;���x�2���z}0������᠜��*e+�e��m��p �I�o,�
��WA�:F96�g��|�J�Cf >�_���\�ZW�늽�� R�2��g����E�A3H���F��X+�'��t�0q���S��������Qۨ,����?���,З�m���U�B̒hh7��	���.�b����%1��J��NM%68 �8yx�1��v�u���e�/i�  � ���S[�^rC|�QW�~!:5ǋ`xi���]���P�ƛ�!������ɽW;�801T�'X�Y��	�����` %�z�(������\G'��R��?TIs���OX����Έ�I^��#]�oVq�\ii�{s)��JK,BE�m�Kg9��懨P��\�?�h[���6?n��.��.@8��[�0��Cf]�M��^�]��܎Ū�g�\0�6����������GД��	P�`33�-F⻼8(  :V�3_,�V���iܬ��[��n@bX��U٬��p�&�a58o����6��O�k��z	��ȟh:���,9I1�����%�8�싉b:^oAQ�ؤ#�{����yb����53�]�Pw#��;�O����YT~XlxVHYEB    a71a    2270(��i=� L����1�����7y�G�ؠЩ�ך���k����դ(̌� ��Β[���jl����ah�����~k���}���\����mv%U!U�����Sù´X��@�d����p��)�{��'�I�H�
�[���|P�y�qJ�9�0k�8�@G����C%�.�4�m�z;���6=��@gi�H����I�
/����8!�S���X�h.�W�N���{�Z�)����lmư�0����Po��:3K�y���,�ƀ|�8x�l���~��|�3�^���n%K��LsҮ!�_���(��D�c$'��C��������SWW����t 1��髰߽g����~q�X�
|n��f�IϜfs춗b y����x�?t$�?xA�Ra�~B��Tv���){,�1��78�����u�3U��X��-�~J!&^&����	e���%T�8�th��\R�3)���Cbag�a
���EC~���1�\F�I��0�	xt&��n#�:N���Q�J���]!�� 2f2���_�Jc�v�B�����w	���ޫj�y%Uq抭��2D��(~*��D+ۥU��h9�?3U3�/�H�z��`�Ga�Ĝ}���cps��	P�l������TEߙ�"����Q���ui� ����"��H� A�3%��@�'��|��*T�o��?L�që�h��?��
��粇��J�k�%�>0h?��R�|��>Ŭ�W��%��fn���|-3�U����!����t�Mw�Jv����	�M�y?6/'��	�����5��q�uPo�(.�7������d ��ŋ�oB+�e�=����9z��	�5�߮�>�0�x6��Kw}X��{Ϩ1�[�l)������Q��
�Ai)�@�Y��5g ~��>�*�u��L�q��U^�D�8�O��O%�ZR�n��@���=t�iD0��2¤�:JZdz��4����\�%Gv�/f��xI#2X����+��WkR�iS1k��z`��1�i��}���j����
�!袀:���B�`��8}�ߩ�����e{�|��3ȯ
��|��pݎNuD�����[���?��:?(x�v�J%9-`{��OE|l� #�M��3.>F�n��y��"��r\[Qph3��FC ���JՊd��g�j�k)F0�B�����E.%�o�v*��k��k&8�K��S�Ht
w�2�*�l�a&rE��R�ء;���Y�>	McK髖,bMP����yVr��H�o7��XUYd���-S�pW�B�6��w{�j�y���
���M�(@I�Y&��e�;���z_hK�/}30�=&�� �n��_��7��E�˝�*/���z���=�G��)�=���D��	R�0�_�260j�_� �s�v�h�%ء���&~���.�u�ш�{mg�,�v���8 �Exk�g� ��K�9��!>�����:����"�h�M�:Ξ� �X�N�l��Lz!-��,U�Hğ~^��\�G��3hס�̰
���|RI_ʜ�;ei�q�+7�`��������$)>*�n���b���D�F��3�iqD���[�o@���OV�H��F��\�9�6�4�l�P7i��}?��7�=����I)�>�o��5��"�gp��*����Ók<x�mX�+�2�wm;tnb�QZ��o�ew߸�8��>c�_y�R�C�]h��x<JU�-��Տ#/_��_��_o]�P�����Dg˾bf��V�]�Fωk*���\P���;v����|O�
+E��4"�Fu�۵~�V�"n&�B�S����c��Ś�~���r��=�l��.%����X�`L�ӈ1%�ј�'�B|w<l������H���˴vD`:���7WMv8����I��%�.�ɒ"P�z���]���O>��aM$XV�ؐ����i�$S��D)5�����=?I�]Ҟ)��U���7�O�H=�16�"��J>��/��5�5�S����l�a6#����'65
����v�E�r=r���R��zP���ϐ�-��z0E�۽��P�c�w�,�K;R�ρ>o�f�h������><ǈ$^��](��X?��~K�0�����L�k?I�q� ��q��@Q�\	�<��B PT��p��Z���̻��]SW1�YQϗ�z]|�;2��Ú�{f�sd���fT�t�ŏ�8��~a�#9�ڒ�3�p9��8���Hl㥯\"y �gq�6-nBU�-[\Ŗ�G�46Xr�K��X�Q�	H���+	�n�)�ìH�����hm�Ω�m0g�+�a2�Z\*_�(��ȋ=��������'[�<`��K�=@�3�s����7"�X}2�1芷�P��N�"_�t�E�Tq��$⫀B>��I�m�x�?�'6nFz���'�ևʇ�3�y�(Le�i�̳y�A�j8 ���В�W��YԠ�첮�/��v9�w�b�Q��'|<����wz��\PM��"���r=�M����I�?:��e���x˨*5��t��1O�w�[��1��|w	��+N��g��ے@ ���B+M�So�dGe�<. ���*������' � �-��������3�:�~�Ӟ3�����S�t�\e[�2�����I�M�Yz���2%⃦+av��QT�~��?�C�wN,e�)	��H˶�O��4b��A�Ï��o=?Ɋ�I���q�t���t�[��u?���q� ���o��	�L3�F���y��
�Go���� ��	�o��8f���q�����I�B{�5���}}*H���Lq�F;���@y��Hb7�6��dG1��	���L�z��1Xa��o�Kt�D��n/T�S�_=�qҔ&N_9�#`�����J\��x(��+{��,�i")�?���Nl#ؕ�r��{���E4�lu�_�D�bùs?�\M�Ǐ�Gc4H�ݟ0.�?��0'��B���\L�?HY�mVk�M���{Z���=	�Q�Q��2M:�Hf���]]�E��'.�lgE�~E��:��6����\9�+$�~U]�z��͞�E.��b𺝍�Y�����\���>ؿ��"TC�ѰF&h�'T�_{�\� Z�L�4Uڬ
���9ֳ��9-�6Q��)���"��*/�!C��EYQ�)�ǣ���l!�����T3�$e�Ɔ@�Y	y�v�K��S�
l�]�����%�
M�ʣ���C�'��B�������iL�2�S���D>�?G�{�Qi�$r>��G�c��>��]��2��/4(h�"����~#�*(�;���qw+��X0O����Q��T�����<muC�\L�ճ��;of��m�n�w;OP���w���o�2�4�#�1+IQZo��k�����a^� �ĵ<���ꌥ )��S	�`p:*m��s��������E#���)�����Q��'�ဨFƗxd);�긹-���e�-�ˣ��)�g��}-�������~Y�1z�&-{�t��.��<qj08g��|�)p`�W��p��i�5��g3+����;=q�!�JqhT�����<<��kG\�	žE�ڥ!�H��]�~�~�dj�p}���<ѡ۫���SR�D,j������6����������Tm�Mߥ�V\��)��N�I;����O�i�w֊�ݙ�ԣ2��iKYB:�O�yǘSF�>���F@C��O�?��vw��}��#NO¨�����X��5o%���}�/o�d��̟�����,�0C�4.��;�N͉��A.�_������N->T�J`���Bu:��_c�I��]裍S�`s����Q�/e9����Ґz�I�h[��<�=��^`����~l~�{]�S�sƟZ ?,�s�<h�ͻ�)�1��\��p6�e�CHa1��q$W?"Tqգ����2؛�?ୌv�4"eb���
���T��6hq��zF��5�tK��,��J��E}�^+�b�Hdљ��;ڡ�Qo��J��aP[��p�{[^�9���`�A^o���Is�g�I�3c��ܲ���AP��N;3SH��3��qp��L�$���1�Ne���}˽��-�ġ;�i|��"U��ʑN��)RlK\�	�n��1�uK�l��%b���{���W%���z�bɿ����<�!�f�S^�WwaF�2r�"��xā�����W@�g��_�T�j�1Q��YRcm⎝3�~^{�M?�m�]c�v�l�}�N�ju$��-�Z���2��ih�6��;GIK��z<������.w�暄N�G��A�#��e�m�����/h����<$ɜU1 ҁ�.�z��"B���������e�6ĕ�����ƱS�HK��>��N%�K߃+',�����M �?��ƳYmj6�)z){����T�t�$���(w����O��G�дV�A={QhV�$�y�G��i@��`d�z:���u��J�P��w?��_�x��L\�x?U����~�u�Q!+��5�D���ó[q���F��eiC�ω������Ă�o;�t�u������\�K�e�xI䕟PB�{%WwM�с&�*d�Q��9�����B3�"�ǖ�,@w�9.�;F��n��!@��PJ�����(q�:�˧��76۲�֬�QH��(���`�s(���;r��<%�	$-b�r}�fp������4ҩMZEA�o ��U�8�h'�hU8�Q{�fVM+���E�����Y�SY��+u�X=LZO����8R|[rzdLV�Ǵ�:�� њ�V��s'�������~[��k7�"g�~r$�Q&U�u`��[(��9R(���i/\
(4-&k�ҡ��0%��03�DB��pvp���U�,�=mS���qB+qF�2Ã��[�կO�ÞѺQ5�޵c�0S�k۱��k�\�Q��FC�:�ſ#C��͜G�Ш,�H6'\d�'[	�$Z������Og�Gw�t�ט�c�0�
l���2�4攝��vlFÎ������V�_爍%9֪#��4i/���1P�T���{�o>8]v=r--&���K�/�Ua_�u,I�� /M%�;!��	>?R%�[�ݣ憰�u^�+5�gp��޺v�es��0lZu1`��]a�0���GP��� �[gv+�����(_y'e\��%4����
�._yf�_��IŴ��d2C$P��p�5=P*���vp:����l�s���O�7��Ǎ?���6�O�`ݻ2� ��
����n�#�>�j��"��
raA��u�M͂�3��ͰlT��B������S �U&�Z��C�G�(p��s!��	�z�����K��p�.��k�g괹'��Oy|�,�5���a�H}r1Z��,��<�
�pQz����0�!(��ؚ����EN���5G�c��=�����>f��.y�|��ES���G�+k���d@��I?f3�78�T���^�ፚz�.�XA���$e`�F�C�����|_�����m��_�-ZniĘ��U����V��v6�e��O�c��z')��!�_my�X�!�Lʂ#u7WXG.�[� �1��7�d�h(������6�:�WT=zg�7�A�jf6{�'�M��Ï��(�y�h��k=��ol��K��Ϸ>��֧B�KIҔ����>�9�x����ƕ��S>)���H�U�x?Qzi��cw0*ʢs�� ��p
���]�ds4�ϵ�����d�ţ��@v�"�Ik�*֒�
ܴ�5���&�Tv���+՘0k6��=5i���ȳ�U]7&/�3*��ݹI��iC��ܔ����_�bg���>c��n���d�R#�$D��}@A�p-m�f,�q��:�[�´�CA��ͯ|�o�&d3�鄆񥠺�$���Ɇ�UoM��N_��L��ޅ�_�r����q_V�iz>&h#��N<����Х�a��O�K��X|`���G�CZ�4)����pI�d2b*�Q��ڰÖ�I���G$H�%� �;y9~�p��ea�C��ɏ�Q�ۉ+J��^�~��݅�e�Y�8'ʍ�dl��S&�V�r�7��yxm�|�Q?���?�ǆOC��x����A�(��xo�q�{P虔���Ѝ�]�F��"��0��O�L��`d�ypC�װam�B��f5�%��ZBSp�1x{�]{��PR8����6�� S��Ѷ/�X�pbP�5�վKZѭn��Ɨ��a���M�0��� ��K��=�~o����p|�ώT��Q_��$��$2�C��)���~��yD�<g�^���>�*ܣkf�匳��P���,��ͻ�h�5��q���ؿچ� ����(�{��M�J|Y(5�;n�Y���:! �G�C��Š�3
���1�|��|�TܻU <3�an��~ͯ��dd��Ó��Zq�`���([C����?^t̔��j�
=H<�]�Q6�	�0-Zg<�α� OOꔏ���a3 ���Ha���@?~�#�aqӤB��;/�о���^^�3�3(o��w8�4Rx����A�-q.*\�d8�;�ov�ѧ��q���򘀷2�|!�q��0��v���7�L֫�	ʥ`�N��a�1��n��8�p�+����'a=�� �����% �z�\��hu���@y��d�F_�Q��D����W2����[7gs8����>�n���{\�Ԁ ~Z��
���π�O,�	��AD厩�4����"��=�����=�2�]�O˧F�JcUx�2ݯ>�^�$�M����iu�U�^K'%d����65��_�!����^�����]��� ���܊u`��P��� ���!��m5$ׄ�r������=�t6��$�_%�2���	�i�dC�T�-~S�N܋GY����D��C�����m���������0[F��?Oα6(�Oс2�[�LszК%rM��n�F9�/`aGIuG�x!��������^�+n�/g�S2�^�"�<�𣖒L��(�ʂC�?����n��@�����<��侼� ��0y}� �^�\7����kf�%AíŘ��n[�G^�E��|�ꂜΏ�@�**���Ȧ�%���k��9�݀�e7��R?�e�q5�[54}!)��w{$�ځ~�k^��`�nTiT����QFo(;l�6_ok�22�"*��h���������2�꡺�-� Ǒ��Q-�M��.[��*%�8��g�|�^�S<P�fC,����4�3���p%�t�5^���Փ��A��FrX��F����RJV ��'N7��l%B�I%a.��b�'�8�aO�k���gj�b�"�z��^���@��^��b���1�!��ϒ���0��U�M��*գ��d[
.���*�o>��f �8��!�C��Ï�ҕŘ����d�>������T�S`$N$�Rptr
��m j�����O|j�p34�ZO����d)�@H�k)פB�r{��z�鰾E]U�)�"P�j�"�,M,��B��.��@��O�?�-1n(SF�-:��A%����V �G�*i����ӫơ��\[��Z[��^�os��*s�����ic�q ���,8dO-�?۾4�\�h҉�{)�5�b��!�D�S�I��<'��NuQbj��}��E�N�Q�;]��BH�Y��lY�Jy���������E�� X�c�yU�c¦H�h��Q#|�f�Ƶ�o	���i�մ�\7�9~�R�C�u�7 �ᵙ#���Q�eKY�d�z����L>�b%4�ى������$w{�/6�ؚ�z6BZ"U��^�w$�Nzc;3,և~G ��=񤻌ǿ� ��-#n7����#�y�k���GY���fփ����"`b]/��qU�`�7�'^�+�P!f��hXਗ̜7fC[J�)ۚ<�?��VF��[���Y!r�j_�%lߙr��uJ�g���U!�=��s(��".�@��5e�<��pL$t��^�f��)'��z��|8+���������r�����l�x���Ec���8<�����0g
9@�Q�d?�A�I�!��ù�5����:�nnZ2���v�&p��L�-�d`�j�.;SD�$���x��웬+P��υ�<4a�12�[K<L���� Z35�0�<��B�����!��l2�F3���'gT��čˍ35F���VI!Z݋Q�n�5	3��b��;�:,]��a��wKO/j
o��^��ަ�S���%]q���^�r���f?4��^��� �K|���"2u�Yܸ�(���7zX#���y"��Ï�'C��}
�a�/X���NU�l��1En�p� ,�)g��œ�T��Υ�^�m*�.��7��M�bm\p�
$s#Ǒ�����o��U��߉����%��\zb��w�JOG�"�P�<���}\@�I�vf�CT�*��EC�I/�4��
���F�k�o�}�)Fp�8�0a�B��a)"b�D����"�瀋����e��	ݨ�;��w륵�Sю��7j��j)�j�ݪ��2-|(O�X��}�C�����4Ro��b�
Bf��8ȫp����0ޏw{�F�+	yy�Q֤��B�z�J�\�6����|6�髀��{�z��s�6�/2�����槣G_�