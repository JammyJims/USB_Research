XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Oe${�W�W?-�� ��^�����[Z���qx�����NP�����X�����}�����1����9��O��n>�
�r��d�<�)ۨ4L�$ܫ����CjzW�O�4�cl����� �������2�+kq�G^}Vw�o��h�\4�\��%A��~�2�]E��eN��}RD��B�í[���(�R�rR�f��N�,��86� �D�e$'ŔJ���H{ŀ�/����	��q��  �w� q&׊��e%E���š�ӂ��M�`l��'N]Q���zH�Rj�	��>]Ը���;�����ʨM�tC�?[�Q�Q#�B�����_|jSC�H:[�1�#5AA�̛/J� ��Z����CN�I�C�^��8A���G�[Υ�"+�+"�� ��v%��r+ֲ�G�q욖����7K�r��H9��|�C���&�s�K���Ѯ���`K���w�~7}�H([ �d��q\�ta6,�c&܎$����V��7:���`I,p	��N��WE׫��ș��A�E�p&#�iOQmJavXW��R,�Z�q��nmN��	���Z������7�������6�?��l��.w�|�z���Rk�!�����]��
��G?��#�Z}�H�>E�������L�_������^o\o��x򇺹�m&���1���|:��}P���]x�|[��R�-k�d�*�>tƂ�B���=3R�w�}.{��&E�D�Y@�\�1��xqt8J
��Eȩ�6���N �M�XlxVHYEB     c3b     5f0�
w拒����TO��&����/��p�[z�c��'{�sF�E�f���t��Զ$j�wRn�r]���1(5�F�a�4/�$yb��0%��ǝ׈)70�Gj��>
��s�<"��+�V�Ű�ǣ�4�2M 7��No{B:�dNk�&��PFj3`h>�;�7F��8���K�5)���5���G��%)�M���J5��oF�q�wq��m��R_?b����y���x6�_@j�	�m�N�i��!��~�SA��yHu0{�XW�dn��l�}|��ޠ'�w�14m�6��wď8Ϗbk�\�~�4 �Od�/����xl��1M�U��~��^������K�Ow(�`Z�;>ZGKG�RC�^4h�����A��A�Ͳ�9��sH���`[��.a�t}reѓ������t��'��ZЌiHjCc���&0���hnyV��I]�a%�h$��ړy�g��윊w�����ވ"�*�CE?8������[����bT��UTM�A�����H���y���+��ď'��o�%��?����F���%m���T�I�����FK}���8�8�'��� ������[Eϲ>�7$�Z��Kq�Z�'��[ڪw/�s"P�k���R��;q���>�x�ݰX����I��?M;�>)�Ϙ���f�-B��YVn��V�Ķ��B֐>��ɰ2�������T�B� 9�-f��H5Z\R(�~"Z.�}�9#�w9�`s�qoq�rz�,�M���@���V��YE�fB�����(��՛����j��Z��©�Z��
#�O|����1���ϭ���K����G���~3��0Z�﷒�������J̤4˕@�w9�e}R���k.��N�>��	��d��BQ�*O���N&Q��!.�Fd�m_�䌋XBN��UC�
�.�&��z��j_lV��j �e��.�|�#h��c8�'�C�1/,���e��{�/V�#�?�ܕ�q�+�7�3�l��H(>���f�ߡ^�cz>AA)��/������ߚl�
��\*���v&�OC��T�YVph@E�"��z�C��1`��6�x�H!~���Z���]��*�o��c�%��7Y��_" ��P��t���b��ݯ
:��~!�m�(�ѷ���2(=+�O��U��P�5��y�?�@�u<oo�e���k��N���	�z�Vz&/��a���:�4�5F9�O+�����;.�>�y�e��%x�ovvQ��$���k����Z�_MW�'~h���������H�Ng���O(�,!0q@z�0�����#DPZ���ۜ�¿kH�g������H&Aن*d���Y֖�Xx؇��B�T�dX����wek�$��lw],oIlNP���KH������347��k_�E2�������>t٤���e5��k b��x��hfc��	v���L���Tx��B�f:��hݱ�Y�re�s�Q�:Dn@��;/�?]R e