XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T�Z���T�а��J�f�!-T���':��v��	3
٦�l�/��Dm�nm lƁ��� N%d�X}}�	Ry�O
�0t��)����ij-g�U���>U��P�X�����x`�#W�*
���G�[E�}}-�)K�o�>��� f���4<��Uqq���^ly�����6�<�R~�eZ��J
=�����c�~�WV�����������Y9�ɓ5'�ѳ�tㄮpǢ�=�t4�8Ȁ22G����1�Ʃ4�|TZ����p���^�ٙe��3� �&p�b�/�- �]�N���)1�Jgzs����O*k?�5��RM�bA<�-���a�p���dwhp!L��\�;A��Km@�0�F��l�����%3�,	�D$�ɇ+�|.iM!���c �]�PG��X�"���?���➝8�y���_��#
�j=��$����1�U�\��Z^J"�BBjZu��T���E��1��R�<���T�z��d��P���G���!*�VH7�?硄X�+!F!�� ��8��<	r��A��C�W����>�/Dg��6׈�<�����秡����3�����h��C~�U���G?�su�w���g*�M'�#{��t��CW]����IX�����C$ik����YANC�'���>�٢�i2lx4�G�[Ty�3|1>A���'�ܚ���$Kc�VR��o3�εC7^4K*��"�ێ�_��VV�O��/���x[�A&��oͮQAC7�}gXlxVHYEB    b2ab    19a0Թ��+����,E�.����/�*��N�������+������CTH�{_B /rǱ���`�Z�C�!����6�d��q.�HOy��B���������w.M�@�i��z�7Uڟ{QP�
����	�cnm��8y�{�1�L<8��e������y���Ӌ�����S�w �1`�	��}R<��b4��O,%��d)K{��W�^�K$�i�i�{d}_��!v�K��nff-;���لp�(��v,I�[���	Lj�x�vh���� ���W7�[ӫD��}|I�`�����ع���ڊy����e�͹<;����oZ&|�
i�W�E!�T��F��N��B�q0��(�иq?S�XkZ6a�8�x+����F '��h{�"��t
>I�1K���4Wb{�ҐQ��ZG�Ί��/PwE{C��7��b��w�X������	��hF�6
!��9�b�&�����L�
/2S�/q���Y� �OWv�_{jNƢ+��׀:7k&�?�:9˟���p�������{�c[��eN����������+{u9���i �]�:�zG�;Z�p���(�	-j�3�i-��������;��� }�����~&5���C�>��G���o{PǢ�b��7��;� �'���$�h�ɥ��gxe @GTٮ��(d�	/ŝc�^A[D=8XA�Ѹ#��֏��^��o��p�{��Y��Y�m�iܷ�
A�\!�Оq���LSo��}�7V�B���GE'8�1hO�n����݃<��g�l���_	�b�$���o��N�l�;'���2��!��$�k�ck�
�������^@9�S����k=A��:$՚�4��^,�@F�]���S	�k��?�0b��3��T��w���U_�#z��Y���d��E��0���u#bh�w:�߮`�Ǖ��F蒂�,�[�F�?��8�7:_{})~�l�0yO^D��5)��E>��j��+>Y��=��@i��L|��_�z�r㖴�ѭh��o4������캼_��`6
�_����Y��L�b�%g�G�]&AߌtS<�̘�~T�n�Z!%C�U5<�'��gp�@E�7Y�D�� S&�٪&���*J��O���E�.Z�ILn4��B0bI]0D^�%b�*F^�1>�ܱ�dŕQ�<�7�� m�����k�\�x�1%'�������8iA�`��rx��W�<��6s�̧�~%��М:�Ǘ(q��g�����'F�4t�A�����F2�����(%�sl�`��W��;�
%��k=����3�Gl���⻱���%r����/W���.�	�kl�Q|>��fUj�1���K�_�\vP�0��C�";���Y跖��% q���Ü�B�ov�A�� �sQ��hoz�������� ����|_d�
��٩�ݱ��J�:��z�>�ۦKaMǔ������ ����M�$IU�q�Ҳ{k�
�!eO�y��5[E��_�`� H:
\*/R�sZ���T?E����S=����9E/R\����G6���J��T2�=��8���&ޱ.�S�
��(!B��(0	��C{�i#�C|��ȼj��$29Ek��J/���͊e�n��/�����6��!��̀�HhS7�� Q���:��r���f4 ���_7UpI[����pB�&au�W�EЏ�䤉��C�9�c�婂�-`Ĉt%�R�_�U��������_~$��3b�YL�ay3�T�`�dL���F�3h���Z��ۚ���xjE����ʡțt�p�EF���Jț5f����u?2����f�z�K�HkE+��]�JȜ��ep3�j�T��hzl�~�v��!��G��@�w����:�đ�5��Fk��]@��;@́Sv�(�Y��%���������۴��i�?���� ~���/5��z
�Y��@O?����BY	���
�3g����y^wX�%�L��^�s�
���k�)̒�4���9�������&�N���1hm.�*�.��J����Y��(q��٘�{�+�4��b��26�D1�<�����޲d~�/Z�G��l"��Q���ۺ��"4�k�0�T8�u�x]I��$�%Ube���k�HE:$�m�{�~��٠��{P�����-A�me����~Y�-�d+^��+���!��i��ǜ�`^�֣^"fnq�F���b�C����o�2#�����u����ړm<���D5���Ui���jVp:v`������r�m芿��^�� �(R������ܿԒks�a��JѸT�w�DȸM�n0z�7�lW�DId��{��qަW�ݎLF>�\�=��|D��$� b���� Y?!�	)���I�����E��v�b�+�%�9��k)/2e�e�&kV-�B�;���O$@CT���`K�9�N���i�A/�����zL��z4���-2�����$,gn�������LA`yW��f7��R-DAPd$��s�.n�Ad�k��TN\>�4K�$�]��`n���v��!x)�h�Sg鵑��/�k4��U�h �p��5{���K-���X�ϲ����z�X�h��7�[.S��6f>��
�~J�	��Jk���{ ´�`�Ge�͹��$l^g��h���n�3Ȏ���u�u�=-����(�|�xh��t���Y@̳< x�ZWK�7aJ,�i�7�Yj.�kt F������Hc�B�v|�_e.��;�r1��۴�ID/��`��sr�4���#��#��Ii��$��{��<cؔ�G�a�s_8~��s������Cjq�"G�D��}��Ţy�����E��NR�Շ8�T���]$�����;�bpxe��k�Q��i�p�d��0�b��$O៻�P��JX�S�4ܯ�&��#Ge4�^��'���o�٦��5�@�T�w�i�UgY�W��3%2l~�㟸�#�����،�f���k���M$GENb�X7���t�r�)�ߗ�B9u&n�+G#�i?4,�[(=s�k>x4�U2�lX�yǂT��Ec�?uJ\f����-�w�

H�nf�Ғh��?�ƥ�b��ٖ�����*dOƜYU#�v�9�Gq�����/C�Bc��&���		�A��J1�Bi�Wڵ�j�;gByT+�;���|��OB[��\���|r��&S��/�4��� �L'�Y{Y�)�sҎ��_w������=��=�NS��弚��Pw�^x>_9��:3ښ�����>���C�;�!����ҜQ�%,��χz�k��l��(��ʥ���5���T����k����Lц�gJ"Ƚ$��i� ����N��8ӻ�F�6`g�O��8�r���1]��� Ԓ��{et�UP>��y*Y�u��٫�8�$��`8�ùS+�
3eޑ@SSˮ�1pz+9�[ ���|:�x�_ؿR�,(m�M!��u�9N.�;Q�M#2@;�9��]�ȷ���~�F56�r)�$��Q��b�5�K����05V���8�c,�͡���Ɲ��n�(�:4���5�bE�2z�=�Őa(w�î���
�����d����`�{�u���c0:](� �
1^0�U�0���W��C�ɣ��3������i���o@ʅ�Id,7�y�㋵�kIe֣7�?1�Ʌ�_�pB��D.\1�i�����i9��U	K��������#!O�&\)g��1�;��`��� o�eiy�o����ʁF;��KF��uA�A�f�S(3�~��
c�׫lk��nȃo��4�	��9NF,*�������؈k"��Z���H�+O��\����)����Z���oj�2���݅�X�ˠ�;&�(޲�'7���;���K$]��]M�ڈ�r?���/�^[�(��a�	]l���;k����+V�f���Vc��.w�2.e��3���h+c1$F_]�|�H�$��X��[��2�FОtG �a�����rM[��N�tf`�S3�z3�P�fT
ݐ5t����]6���CU�S>EV��Gu��み�x
Vr�"6� �/`k�.9"�$A��--�ԅ��,��$ŭ��:����� ��$7t��$�м!��5?z�:��d
B�1�ȫHa5yi��~�#;�RP��$����iz�2�c,�|�������Ü��sҮ��������e���Zܰ��x���t %�����;�vUuX)����A2�'����d݌I��Tu� sa���Jx��eS��:5�LEl�>h�[{oPS%5F
A�{Gv�f��@�*��݀�+N�?L?�g���   O��[79w>G��G���w1���DA�e�Ύ��!�H�ʛ���|Xޙ�)�h[z���{!E�h�y>�9rr���6���P�L���� ��;�qE��O�v����H��kű�2�,�>�Nsu�8؂5�g^)�1���'ciK�'?N8��$��\5��f���FQ��t���N��J�M��0x@�9]��#k���}�x��G&��+��3ҏ���@�����x�
�0�����1"��B�Pˆ�gO�݄f\VKD��
����>��ј7-���1=$��"$0���z�t��<��W9�Y�3|{�R�&�h9ز�\��)-Uhn2Vi��{ͅ�n�%h^��02��.M#����G�̵H�"�D=~}�����p��!�.��Ԛ�X~�2��o���`��6��n7+a��vٗ:f�P�X9Ȳ�piO\��n��]�	> �k	��te�$�����Y�	!�`'&������[����=[�`|.�4,4V(j�ܧ-�����I��& ����K�B��Ըۛ���12���w��[RK%�NØ]F@�b��a����9׎�`�V�M���A��Ҍ]} �T�~�ҍ5� S����Jd�סe�=��M�Q�Ph�����p�d�U�����U"�����b^���ob�:*Aw74�]+ڽ��P�>-=0�s;c��4{oj�i��k}��d��G�,�"m<���Y��Z�_R>F2[�b8���l�31p�E�Z��ŷ�'U�e�&�L/秹aC1�.St~��C�$.���W��) ��8�5��$oI�W}yy�kw��@�v��Uق��(��y�xT�ME��8��<+M��*�	��X7!r �j}r�|�ۤI�:w�?��ۑBd�u�:�8��A���~"��)�;�n���J��J�����x%(��bL�`;uMn��w�?i7Yr\�ȼ�
��k�_���^I���2���3q��!7wHB�2E}ݪ�������S��M�Iou��<�=�2u�����tHJ*&��d�1����V� l�w~�6�T%�v8o[ h�A�=䶠c��{IGI6��,
�N��a��"l�ܨ�j�X��;�jK��3�+.�v��<6�ןpڎ��|���x^1V��/��&݅�8��7��㑱��1HCp:�M��=����Lx���P`n���Z�x�C��������N6��CL}ۛ?v-� Z(B��������s5�<�<��\
9�|� �[3�:�,G!���# z_G��Su�\ �T�Q�S�e.���m�?�*!�6&��z�Q��#P�����a�Lz*�G^+eȨ�3��f|�ߠ}~�:k��������*::-������$"]8Tb ��e�%#۟���B'Ƙ����gC�p�E���$ad34�����y*�I?����cf;V�ϻ��9�{sS�#9r+��X9	w��7��{ ��H��"�c���>�TA�CbQr���oU�n�XԴiy������ȟ3P�@����"ݷ ZI��� 0���MF-
T�@z$/����|{T,�IW��o���~������g�a���?�Y�j�(n�$��s�ʂ��f&�Q<s�t���3.�W��!87ēt��J������G��n����i�k�.�d�b}���̓���X�<9֠�����yJ'
Aot���~ѩ�oi���H3?�`�r�b���Y�8ٴ-�(�O�OÐ�����gȆ�B�ҧI�C�j��Vun�+յܽj;����uܬb5N�*��xRm�{��Op���7�0B�ڗ�.�1�e��j�L@9�F`��Q�42�#�Eq.��L[f����X1����1����Ug��ZFӮF�F�jQ�4)�_�o�}��״�(���?.�%�㴭}U��Ӧ4K4!��N�e�$�C�xc�wX@��K�8$�@ļ�Im�2`Y���F*S� �eK"�&u��b��� �l����Ry��F[V�Q�'��WS��^��&�߄��%�����֫�����&L���<���D�i�����oԍ�M�=��C$��C����_��&���)��p���-�Q�mUV�o�e�<�OkV����8��_�8���#��j���m��Ms����; N�V�c���-b���^