XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���4�y��=�V��z�=��4y�E`ݮ�t��8h�rf9�)D�j{&�wB7ǴL�xp�D��6C���h
ќa�f�C�%� �W��(��f����L%�P`j���9I�-~�����_�Bvv������SD���~�����7�|P�AB(X�����c�'1�5*#�rSID;!m����ۄn��/=��KS�j�z�@�U��Km:��}e���zN�,mc��P�6���~��S\��s��	��M�w��1K�)�*#�?��y�/�1/\��,m����|�!�����A��S��{�`F�4�6����fm7�c�wS����S�VL�A��@�)�x�x<g��ڏ%���(,Y�e������n2,��ݦoh���"`�3��)�R
�/���!]�]��� b�XL��G�m�,�p�̏V'őB{
���=w)QdME�<F���oi�B��I�Z�?_��[�i�	g�槇H0�ˠ$|*d� RU˺����|��"�ʎsP�2o?�߱찇1���t��Ff�
��$����
�B����.��AC�$��ृ>���]V�����_��퐵�A0��ҫ�猛�̴��k�A���o�|o�^����d���c-ܰ�>�r����֧��Lp�?�gCg��
C�!#�UO�0D��^�����t/2;4�͛�b���[���c�3�7���^����7^��2}^SZӹ�M���߄O�>@��5Z�������5{�k�r~�q�z�WvWU�p�eXlxVHYEB    47eb    1000��A�Rf����y�vr>�kJ��* Y���;d���3_����������m�SN�9 a�7y?��5߲=�#~��:�xp�0�����9�:8��Ź��"8��hC��bG @5�K������~�P��:��&�΋CT�����yEK�������sT�)sf?|f+�a���=�ª���V�Cz���k���EK6#ֶa�v�H�DHse�[ɳ*|��L���N��D�<l9��L./Hpa��>�U睗�s�h��oA��̌�ԦOO�^����w��1N��]D�z�v�����5q��Mi���(��0���������p��j���R�T:;��d�@��~|du/-UB��$���(9�8��r��V(8C�?�_�r>
l����U'�@�r8��<�ߚ���/�%�F��=��t���Wԇ�c̚�f5����Fw�ϡ�^�Gz��'j��_�J�P[`pۭ�o�P�������X��F����E\`*Ƞ���FR�?�6�3Pp��J�?��%�_�l����
�􍤠���Q���|7<+���3s]y���rɲ�7�j�*�ȏ���%�߂���҂����@/���5��kv܏�y� v��S��,��f�\O��E�d��jw�@�(���8������6Pp !}�^	E��	|H;�dQ�#F{kbQ}���1��E��,eͺ$^��\ǝBY�X�U�ю�������pֽ���q�'��I���v�!V\&�:�+�>�!=_�<n�Ts!�
�O�Wh�-���b��*�gZɩ����D�xD?*�n�}*n�~�y5(�zlIlZ/믋Y���'�	�8���o3
ӂ{DAE��-�"����� 1'J�ij�I���#��N�j<��W|�f$���d��k����cm��>5�C�(�	E��97P���n+��g��5��x��y0h�k��׼��h�e �#��$DkfI�vt�SO��O|/"��mnH3f����%͐ZS!����4�߷�Y�>�� 3�S�/�O�ۤ�R+��NZӣ�U+!���K�?��|��k��j!"J; e��λBd�$m��1IO�H��LSS���Zl����7'0�D�wV,���9�}:?9�K;��Z�?�Kc�N��t�`�"�\��K�Y���G����<�����}V�(tRPa�%����*���s�)>��g�ɓ@� oD �]�o��G����T-�0gO��I�;�/��#B���(g�O)0Q�z0�oo�A�r�Z�攀�m�o�����Áx��޻M�m�c_
�۔���*:�(6�ۿc_o)�̑��4;�?5�0�n:�j�-���ٺۘ����6�0O`����A�ҔQ.5,�'ڰ�=.J"��
ւ�,�X���
��PMx���!�}���6l�u��j.#���1��0c�Y$��*�Zs�+T�H���3��"u��%��-� z{�n�#�QJ����b,�[��'�,�`����/1(ѝ�ǁ 6IHY-�DUa����MAV������ ���Y�9C�cά��o���C6��	,t��O��q�ؠ�:4�Jo�TG����wʕCJ��k@Y:Z�T�G3��!pSh�*424� �!D�����}fk���\.������_�Y�%�Xg�4Y�Sc_^fVD���q2G����|.�0���k�+'�������j'��VR3�F�~�h��+��T��o�on�7֞Xݻ��Bp��M�j=( ׼��R?F�^j��zeK¿���{�O��=����1�B�PF�6�B�&5��7���,�_��8צ�A�j����b7dp��]s��� �)�<��۳q<�����R�m���rT1ɱw��AP��J��a�/Ν3>X���._ʓQ���3��_8MS����J��|#&�IqXbK�RgێG����B�dŢ�9Ɲi�Ysf�����H�YJqq��Q����!��$-t��mp �Uϟ<"�!r�I�s��(�H�W�������n�	��Fd ��N�:B
xW�����D�%sK�\�J�Tա����?�`O�́�Ǩ���s�Yԇ���׵�C(+�m��޼M��7a(0�NPc�5	@	rm�X����o��e�e�E�]��w�I���"���8,���99���Z���..��Y�?3����a��E�~�b�e�A~�!T���Y��k�K�s�чlJ�N4��n�ғ�@�*񏩾��EG����?
w��{�Հ�!TL&�+` ����,���$�@Ϭ�T�I�(�iT�����<[��դ�x�¥ �fsM�1�ļ_v��2."�"��R�3mv�U\fs'��/�m
\{!���w#��r}��;k`Hxlӣ���/�"��SX�/�Đ^?fx�f쾐,*��(e���D�_f:G9��eM9��F���mv[��L���ن�Hܽ}����2J���Mk��ͨ3u��M`�:���r�
t��Y�����N* ֨����P�4x�K.��@�:G6��-�v��6��\��P\I�Չr���d2'o����v�_e�L���FR|����f���<��юG�oзd���z1A184�M��84��J��Z5N��&��P���J���Ymy����[�β�L��@\y0Mא�� �F�"�[��=8�-Ei�]��?l/BB^Zg���s5��[x	�M˰���7�c�_����b,.�~a��`�U�����-�B���'�b���QFg�o��uM/��Mu��x�D�;ss�n��;ᱍL�i�0 ?���2���cߢ������s|؃�Z����UK�U���[B�n�BO*2lS�:���%Ah	�[P���=)hp�[�\pdZzOLh"���.@��;ꩨF
�e�X�c��w�5�B��پ���&���+?��)���8e���OB�jsb⠖W�O�d�K������M6ٛC^�XIwᒆRB��b�-�i�B�ck�U7�H(�o'���	��#x~g���U�St^��R����l<%s6�`TI��`T��6.|9��Rb��a��}k�p�m�����T�����1:��r��z����V"b�9K�0��?|�Rx�6��`�9"�h}��^�!'wD���d���V���|jT~D��K��
���n+����0�N�:_����=�T�Z1�kyV�*俠IbF��7QH]:g �&�,R�Nf��ı�̽rc�C�2Dpڞqj#���W.��ha���v� bxZϬ�O��|{�I��c�koL�*��cD��3�"-���稉��[�B����/k���<�}�[��!LS�#K�F��A�=[�SqCSaJ5��N��ۤED��jEN&�ľ)��~`"�[_���+]���l<.��=�!M��Sr�ib2�����XҬCPDR28eKgi)Ǽ�-*�αEY-���� %bک�� -��ơ��C$�!�<Y�\����?i����[q�H�<x+����>EN~���}�Ee�h� ��O׺�ћ�j��G͛�V�(�ù�=��󨛡��0p*x(����ON��3�`��mÛ�A��w���!�[?�4�r#�ڈ�:���ж��-�63��_��{��b�%}2�*�6�@��k	��FT�x(�S手ffۥ�ZE=�2�ҺQ�8�7i��y��a���>��ǩ�1���������r�č|��6Ьb�r|�X�hR�5&W��ՙ��Q�M�g�
]9{���᠋��B��)���0��Bz&�,����f���0¹dK�ֻ�}�5C���Y�h����Q��S��k����G�������;f{��)~�\c{? �$�̳�h9��Qi�3����M�s{��LSψ��y�m���I�,�VW�kOKGTwT- ]������:���=A!j:�&'j�iC�H�gr
Gל�Bz��W�H,8X�� ��ਡ���[.iF6�������bņQ�ዳT�6_����&9������`��Ʀ��2�N�