XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G����e�K�[3��͍z,��B�O�|����8����V�]��DC��'�^i����8������FA�C{�՟\r�}�S��10{v}0O�o�uy(�4�>N�	���a/حL`GHCh}n1��!�Xk�x�" +�G+L��	�'��o����!~Gb��=���l�7b�CPC�u�0�A��WGh���G�������8����D5m�ʞ���|`_�Dr���*��slMY*>��;*�[~�~A��+�'Gڲ�ѧ�C�=g�[8��UEB��V�>Pګ�R�"�	��Z�~�&�xs�R���7�V*lUx�N�v����(O>�KФ�������j� �1�0����E�®��d�ܳyu���?/�˔����jC�[�6Y�y���oKIO�����F���C?w����yXX�q��l�38��e�� t�sj�A�`l�UV���l��Lwt}�" e����	<}�o~����&`V�I#�;w��.a:�Ƭ�&=���1��j�!�s�: �"�+ؼ�����U�̣���J�%�s��(yG|Q���TLJq��[=:�@��nP��l:�r�~�Jo�4�Y(�2�(d!T��/-��:�^XZT���#O:�?-C����R3��u�B��~�|�+t�!	�m}��k��y��)=g��sz.��@Ǒ�Jz��n�f�+
+���6�gly�z�uK�l���.���cQZ�I��H��b?_�m��T����XlxVHYEB    f4a7    2f90�oOH:!t�&��DHg]�fG�9D�����ҭ���"�w6>�<(����u����.L�}#Kv���bm�{z�.}��{��f8�!��6[@�s`�W4����,(>h��q�`�h�s��r?&tMN}�h�Hk�$�ah#F�o� Q���[mīN(^�HU�er�h�-	��B��rV.Kj��~�����Q��Z�l�3�i�
�XP)3ԝc�~�Qu�E�����ҳd����hQ�۪?Ƌ���x?����b�p��G+j:�ơU��׀��#d�	�����s�KទQ���V�0[i|��*�
R,{���%�"���_��|-!�>��A=e�o-bŕ���jLM����j��8P�(��$���9	%����2�z{q'�a%�aG	g���朗���
=�Z��F��Ͼ�Z;�G!P��^W���T9GE�(t*hV��� �e�7�g%�կ��L�O�_�Ca�]�x`��|B<�g�TH�z�f��e�u� R��!���$o��%����V�IYPW����!�<'�,X�}"Y����9f�d����VΉ:��⌵1�B�����?E�˩�|5�HE��9���u� n��!�1�N��<OgV�XB��4��=~��E��C D�r�FۖG���-A�ʏ��bL�!�Z"u���i�����������X����;���Ԫ�i:-EJ�����!����r� [j��Ln\�
��?v>��4�%N�1�.-�+8���
̇y?�Ij����s����Ur��Uډ�=�v���
�)�&���#���=$�C,�\�݈��\u�M4��`X����%�qc�37�Qk7�T�7��;\��X�G��MBّ�o^c���%��ŸG�K�2�q,�Sd;m$(}�����t��٭-�!�S��T�z�YGs��)T]�/xH�V��Qx�e�y��G��Hǖ+�z�O��ϬS��)���$N�i��;y�
�ɍ^sYPb�YhU���v@�Iʣ�����
�AS���`)`]�J6�R����T.¤/kR x�}�b߰���*x��F�w�eBU:��e��%��cX��B�Ȉ�*���G���<��.0z�U\�{����2���4r�F{DS���[V�fV\-@!O�ӰU�Ă�P���L�}�U��] ��`|J�М��}��<pHƜ�&5n�'FE/��}��Qσr/�Q��+�H�o�^`�@�����ùs�J�o����Ҫ�ik����6�L�p<���+��v�CJ�6	��W�)�|\�T6*�9_�@j\{!��Z��t=B�&�We� ��)�C�/��s"' ����d9��!a�#aUDMK�)\	�%����EP�0B*�$�q�x���<��wv�Oy��޲RMޢz��|��@���0�� �.<�ӹ+���NY7�f�n���MS�i�H���ç&O��h�_G���;�#"�P5�HR���R����yF�|Q��d`�_Go5�Fۺ�A���=�����R7|�;ʺ�kN�ҹU^��U%4F�>?��P����
�dXқب\"8�n����Mk�oʡ�75�^��}��o�;|8��-��� �XVzɓ�`UPBzB9���`V:��v�n�w��q�Q�'\��4kN�+���R75 �͎����*l�vA��[oj)�lFo��eF�i���Ԑ>j�#�?��-z�A,VS'���/$��$~��1];��z���K0jr����1-쁔��qX�����{GsEW�Մ��x�)v����D��yd��lnD��T\���X%j���*!Z�]�n� xD���q�b��m8�k�@��/��=誮"y�FQ%\5���m�pFW�ȦY4[���;#1��?� (j�}bҿ=��������s��.�bK[A=0]��p�␬<�
�R�<m�r�4��S�+���=`�)��cE`����[��M�Q�"lϭ�n7���Uw�Wm��}�<���f�vTR��,��
5^�zp+ul`���T�?w[��\.(�_�̞��P�We���M*G��J���:�q��:�!J%��l?� ����,�Z�����p2��mK��~��f��sV����^�b�/"��.QCc�6�ț�Y�8�wNz�ڿ��\�f����+5x���}�;+�t r�i�<l��8���	��E�px�����;o]�ΞDz�������f��)>���bLqh�~|az��%�1q�����ˣ�)쒎�RR.���h�Rv<�<���Z��?�����~s�]A玞߇e���UW�����a���ML����-�e���-�"���&��(P~��9cu�D�Aox���+QNzWx�^dD��M�#�)����8n���mV&U�<�rJ�\��+��������+^7ݞ��O��7�??�7ԁ�>��?�U���m������Ǭ�o}{q��;�$�)������PyS�WA�~dݐK�XPlO;�x���ʼK(�$D�_)]gKH�(HZ:@��n�;���'�>���K��m��F7Z|%Z���n
U;��,�8�	
�'1 ����V�-�&P/̍ϴ�*��}n�i��+%�7w�-D#l��������C��T���\+�e(�~*�k_���|I�����z��1���*����ծ;mB�苯sY0��\�ڲ�����@y��~"�+��"�����fw��?��޾�#WX�r�@:�FOF�ea���"┢��v{xGrj�&]$��(�!���U�e����X#���R7���5_�C���Rd�W�<�fYDV�u1���h7䑊��/R
�m[޲Lrw��G\}]�z��'$/�W��-�<1�23/���F?�>G�lfV�[1�5C�9H_m����|��tV��C��@;��d�v�R(�1�*PS����Md�'?obԅm'�h���}�ݱ���-qv�����w>�G��3+�o#(�� P��u��QR��j�B՞"���!�E�S�б�����(�d���`�$R�!f��b��;�!)X�Z�ܡ>�����K|�s�U���J­�+��5u������>Y��F���cܹg)��C{�n��顯���qٝ<�%��`3�c
�p7�/۟M*��[6�������&��X)�+�A�� ��OF����{�R��j�R�|���+&>2����}�ثi�vB���@̢H]�s)���Qt�35l��J3��-�L={W��"� dX����+���A+j�oۥ���(g��t�P�� ����q�h��";��f(w' l>}EY�,���9�}$m��/��|!��(`���a�x^�Trջ��d��#9&��W�C�7vC�5� ��f=
���"�lD������"�3~��R>_����\}��\�NJ%a�
�WJ?HS^C�#��n�O�ӈ��U�1�E���}�+vPS)p�s4�Ȍ����n�#,x��?MXp�ֺs��	3d>���s@�s���ϹHD��v�bX"[v!w�?���C'�0o9��M(��p���Ԅ�F,h���0��CP���*TT����̓e4�ݩNЀ����F"�uwOm�$t���Gc�����>v���CX�s�]ѸN�l���Z�V�
f&��;�'6�,��ͦ{�p �?H1����5� �9����\�d�.��4�RDpd6��+�$�t�i���f4��Yg'h�*�/@R$�qwR���r��h����Ժ=�>0ܳ�Ƞ,��P�':D����@*
7;&�΀[���L��4��Μ~�5Fh3>�*8F��/��t�0�<U�������K$���M��``�S�$K�Q�ܳ�jXQh�qf��md��&+J��LQ�����%�@k`���>��[��!EK��������JYX�RI��Z�)f	J�!s�1��D�s'��@�Y�N�ƪ�&j :����-N��S�ζ�>��=�v��|�-��m���L��H婼�$�npv.�T&�䖕w!ȇ�p㜪dV��w�����-��Gw��9��%G�N<��ԂOPv?߰3t��y�16�@�a�ez/��l��Q2-�JI��y/8���`Gc-��fa���;TKnB�cc�F�� � 5Ħ�Y�UJ힦������A]�c�ٿ��ޖfZ Y��,��z�VG>����,�\�F�k���F�VJ��F��\����U�`��7ؕ(����{�}���@���i^}Ŵ �w܄��plFⶮY�k��x�V0��&�;�s	��}���,�j��L6�I�����	�Bi��]$���Ȯ�J�m�0�*�5������5�a���ZK׆�.�J]�n}��Y�l�G��1bg����t[��0��{j�:nx����kF8��㮐�2�8寧*o��x��g�SԌH���,�b�?&<�4ۀ^H�S��b�M	$���3FS���6����������`	9|����MK(��k_Wm�P�*����*����	�<�U�Ԍ���o3��b�ܝ�$�f6"=Z�ĤH�T>�u��.�c5�w|�>J���xS�W3��s� ���wdE�; �o��1�BW�/�BI��GR�
�'�[h�'������$�Z�N�}	�m^�����Ƞ�K�:W���ĬFk�#�J 
�[��*yi���/�źTSS�%�Z�|�� �JrP����vٲK�����&�Z�j��������|���-A@�
�39ϝ}����.}��H?���L6ړ���r��$$��P�׾*�ª�cJ���!Ȏ)b������O�E bf6� L�$�������|��u��77v1��\���o���,L�����p~���wo@��৊+�d=s�D|���]��`gΈ��zS�H���ԥ(����
iTR��ܵ���Д}��O�7iBc�r�씑�������\J��A�:��AF޺�1��ճ��{�o�kY�wb.�-���<��/�A�M�QK<��P���m���;*��Q��:���{��E$^>�`�b��nG�jp��o�8Q�Ϯ�.�(�Q0�;�( 2��U�z�@�Qi�-r<m����d�3{ܐ����j�i2���;�j�zh9>�v�!����j����&�%��UM$W�טUv�c�Hf`�~��Z!��X��L	��)�G�Ԉ}3�w�H5����)Â ��@]�,r�V���8��U/!�Pu5+2mς3�dAϣ�axݍ5�h�{��kM�F1��7�6I�&�;.�>-��� � ^����g�_��x��8�%"���`ʲ��?q��)v��Er�cdm��^{ +GS@�,7bb�x��g-2]�%���9a�iU���='�32���kb�u�%����*�]5L�`��h��6)AA�0T�*�x |�T��j��� y ˴-���p��v)�}�z��Oq�	:����\<8Dr$�6�t�`�4ʲe�^ʴ+RT!�����C�/�-~0���J�9b�i;}iδ�\�~i�o��AΫj�*07�2�{�Y��3�z æԄ�׀n�����-��iB�Wc;��[�ܮK�C�d_�f��x�]]�5�.�nI[�{�^h/�@��lR��;��P
,�h��}�G\1U>�7v�����XJńw�p�H%��L�5#n0�[_w���2����������S���Pg�u{��yt��{�{�]�񄷬����cV���Lb͖��T ������>�E)u��$9"���`��� �|��#��$g_��AT)͊qϿ��NF���� �~n�o�V�7�X����ʡ�"ى��
���ʰE����\�k��A�uP�)�^�,8����J��v��	�_2�e�6�N
��[Е�<M'A�6��R���Q��I�ܱ�Jk*hY��#��Z�uj���"�d��T�١�)`T1�sxB���wU�Y,g�T��Q98���q�	w��ޡ"��D
�M�T|�LX��߷��ӟ�Y��&~�;�:>����������W$��+ ���] 6�'s�e�`�0��,��5r0�.x��.O3���#v��F0��4�wA��a�^�Ie�D.�:�(Kʊ��%�ؿz=��
{�Ϩ�� �8�������a&#���� 󪎙����K\�=�_ŀ�?_3�g�t����2vR:R�G����[�̩���=Ʉ>>�Qk��/��i��
d$��↷�ߤO+�f�m��b�$B{ԭE����6�T�����Ox�z��u���)�y�ӯ�p��������]~��/�JnQ<M���FL<�jҮ�{c�����&����Vlҵd-"d���W>��*'��3�=���:vjt���ŭ=�6�r��Td�>=|�����mq(��xIB���ƾF<�T�
��I�}l�|a?T�����������:R�C.�K\/ ��Rx��o��E訶��ى�~0]�R}�$�N�`�|�[��/^*t�h5�8W���@��Y���;�Ec;q:	)��xB<$(�C�)EdVU�g��F���T ���8v����RȎ�+�v$��M�Av��	�+�Jk�Wa�R::�ޅ&uA��~k��U�T�����~NӬ[��L�b��l7���,�g��FK���82�Ʃ���[5q�������;O��6�7_���ca���1<թ=���̿�K'���@�:9�f|U\���9k"ω��Cn��\�95Z����:Zr�3I��U�eO\�,	Շ9_ܗe?I;�>2��0������.+� �zb�%RU�+��K�@	t�����K�9/ݰL����aer�ӟ�Jg&�u΋�䒝G�2%M�nS��u�j�吪^� C��ٞu�/��BM��E��|�)!����ӑ�5�c\F�Z�55X���h�cTsg ��^��9�Y�-ͥG����S5q�_����#֗5�H@����T�hmJ�����[XB�O�EDF�Gّ��C,4S=V���4wa��c�����6�\}L��ۢ�~4ֈ�zլ��o�NtD���!�����j�n���}V�+ٶ���7�f�� 3T߸J�5���r�����4%�O�����4@��榅Y�/�3)�i_k����ay����JPo1���M�s+�ɬ����QG 2�'B� e?��f�s�;J����'�.���Į�KULt��3��N&�TxN��U�\��Yo�(�^�[�:l������K�7�:���"��=�y��|�Z����
��Z(�2�N��켽��ݢ�? �� �Z��NpjcQ�Si�^��L���z��s�Y3i�\�Jq��"���|3���skF���a�/?1��6�����3��mp0/WuB=`���X*O��tr�,l ���_��6��}�ڻ�!U���K��#T�Šy��)yw�[��\�7�����^��ՙl��k�n&gt8�w��`x�'O<Ȓ�rD���3x�Y�B؍��OiY�Mӫ"���O:Ϩ۟%�km�\?dF�2��j4L��4	�L=ނ�Dj�5(�">X8����8�D��� ����G��nч���,T�=�y$>�#Gq*O�`�J�� ��R+r�g^�T��X�ndT7��>qD�n����g�<�V��[Hd#˯��-˺{�Cyۓ�֜Ja�	n��n�a�$��IX�ժ�3fT	�\RVu�	b�u//�Y!�4f�!q��̝M�q;�g�L7���W�F0I4�߷e�pI�@���?�z��p<�N 5�;�|{�OE_a��]7ð�3��9z�V�tF�fVX����.�_��י)`ɧ�8�`���)�z}��v�b�W:��WǠ)Eh�iLQ�����[�`�-Aa��N���4aC��g��{����)In�D�DY�����xTH����vĥ(G4��ZЍLXL�ԟOJqȭZ1?6��?�K�=�_Lk�2
-F���`�ҭ1��2��Wo�7�Px]l�}$D��t��Ms�;2�{a�Um�J-~Ǆ�5D<�U��-�^��T�R��x�%M��o?�����X̀�j�>C �y%BjzoWN7��3��"x.`k-)J���6V	��ۃ��CA���ȗz�_y�2O�I`���>�7iD�s;ǩp�9��%�d�A	@�r|�qbߥ�)א ���W ��B��%��rV�~|4�s��� Qu"��C�N^�yn2�XL�<��q+�;h���]K�O��FQ��`��``�4D�)��Q���qd�ǲ��z%��6zw�[F"��c��vߋ�m�hk�N�� b$�nz�)
�fh�z]Q��?8��D�C�H&s��s
[��H��c4��ݏ0�����mu�X��W����9���t�*`;�K���Lk}�����8��fE �
�Ǳ� ���N ���`gX[�]�����{F���-onF~�'�'P:��0��z�g���.Sm���zk�?-�!߃��rKt�I�s�o�"�/��H<ڹ)����\�݈�4:��2ܐq_�����1��|�܄��"��L= ��9L��|g��q��9v'��)��`X~ML�#��� �3�%�t�j�#R�rx{�O*$R����h���u�~�D�H�Y�w�}�N��ܟ��ll8��I�Y�͛�k�J��%:gDp+�o�RB޵�����ǃ��aܗF Pݡ�j���u����<��R$�W8
�`� ��ۢ�k35�s��@������ו�#��ݥj'G]@��9�}=F�r�ċ��,�t'�V��E-��]��2����,,�����ۦ7�5���s�����=��f,���!��I�L��X�H��D��Ʈ���=$!��}Hܑ�t�Ҋ���p؇kMk�L��$�'$�S��G�h�m��C�~���$5�����A�Dw��.�@����Y��&�B�a �9Xv�ڼ�Ə7��Сe��9�����e�Ý�I����(�ꖾ䃈�B%�L/�����Z�&YKJ�G�$���/l��N���K�UD~��z�Ұ)� pg�#N7�'5�_��t��}�'�k?��� ���8&��������V�u�n�g��}#RaK�8�e��xW)��w���b��@Hm&�e1|��:�����1}Y[������TO�b��1�j���xh/FGE.y	��7�!1�j�}�2	s�_������ਗIJ���{��"��(�'�BVJn����������|�G<�� eg��W?k���Q����Y{��
�Ro5Z�3��NR���k��`0i�}u��"?խ���a䓧H%�*<���%��^�����F��O�h��[=�+l	�
Mx�<�+���K���4vt[c���u�fZ�-e^�������;���v�U��gL\�����m�$�u[#�V��#^��&��Y�N�ǎ6��3-�>W1j
*��k@�w~92�L�������E�U �YB��V ;\�5��h���?Ɲ�v����\]Hw�GV>��-��ޖr�=O�-�2��қ��T�i∪�D�뤻�-��#i��k�Q�k��#��[������<X��
�v�v/�%.A�5�2�߃ۀ���/>�Hs4�u.�w�di?:=I��Ǉ�����EP�l����]��~����<�C�z�"���~�lN �,�����t�H�fs�l��ô�{Y�����y[��œpkn ^R|�gy�y�Yz���1-ҡ7�Ց�0����z1:]8��V�p�lʟM��*aM>���X�r� �R̰rPO7Z��>q*�L6{�c���U3�VD���{*i���h*��I��e�@�ևu�k՛��N�j[R�`ڗ�`0�/Mn�*ʵ|.>X�������h[�fβm��N�#_`���!t8��(Zkyu��Q���Dě��٩)_�̙Bȗ��4ґ��l,�
<�}�e��@�bbĖ��9�W�A"��<;dZ�������T�5jd�A���R'i��r.}�G̺��ZÙ ��g��b%b��NE98�a�-�����OL���rƋ�zԾ��w��y��l�gTUn����T���h¶,�ô�̀�SuVLB���_���'w�f ��;s��p/M:�`��'l�-��q�ֳU�pċ��_u�bQ��E$i�xu-b�\�u�s��fS����ZY�|\�ΓS�f����I���6�7��r���V[�7�x��[E��@����ز$l�]��;��sBo���s���(Յv���s�����_B[�bHh��pI�3K�[q#�a�v��,�[T��PU�]�i�2%f4D�"c�G�H�s=�8�>[D� �+�B��S����pTn����\H�<�q��濐���|'�g��v0��q�\9>�L�T��j�n֊c}��T���9�׈6ܘ���������ܝZ�M|�p�r����t�c7?�pA�`Ǣ�!��H�У��|z��	�����`Ů�ä��J�-�_2q���ȯ;����^��2�d����n��Ң+N�T�2��6t/�('���'{��CF)�TMf�o��\fA��0O	����vЦ���c��;A�<��$��d ��cӟr��[��C{�j�#S�E�Y�#��`����"	r�r�L�'`�j���e����"P���a�:���D��>o�ʫiG�j�ISc�tA�t��"��n��Q�兪�{/g�#&�O�7���L���w��w� X�&C���.u�~|@Z�Q=�[���3i��e���V;"_��@!S��n�fMLA�&��Q�.��t �{������V�E�Dw��X���Ʃ�~��;I9��R�!<\1r;�Q��83S����Z�72#ٮ��ď4�Έ#�a�y��X�;�us=[e�`��p<s[{�������/a�9��ʒ
B��g��1�6��A)��:Pn��P���pR;�2N�9�%�ڏ��x\��|�JK�����jA��m.q�f�=,�Q��I塠�����m~P���Ƕ>n�w��al�4�F���|����PtP����#�ƞd�׵�U}#o)��K��0y��c�$^��(��vx�e�y�%Wp�O0OX~�	���҈lW�/���Z܀�����X��D,�M�y\�Vڤ,C,D��?�^�[���~�lz V����ir��F44A�Q��7�1(lu���O�+������ќC�"������/s�SHBn#4�����Z0���ź?2�E��h	*�X�*`��d�hK^v�t�|�9*Y�j�r6o/�*�=ҥn�R�V��G���	 Tp.���r������)�6ucFϔ��%�����j����G0�F�YJ���%�}Jۘ6j[j�r;�z�(M
�V#��<�ll�uzYKs|(��8���r��2��{犲1��J�Q�*�$���(&Kc<�G���p�|:�2�T�s��r��q�<�ym~}�{$,;��jt��O+6u���<�5�n/+�{��>���1�[������wǔz8<\�\S]�'�d� q��V*����{q��%���b�uр�Q�s��|����g_.;�Ё炨�ƜiT"��RW�p|��D����=F�ܶ%B��
�s|Ԩ��D�0wOx�@w)!}*8����!�F=�G[ėϣ�!P�Y�t7=�u�8�A �X���}��CЁ����ǾM����o��<6��(1kN��%����lmG���E�Y��%1�����#������A1��%̉j;'Y�K#o��#���ˑ��V6@K	R����?F"R�_��rv����T2���D�2d���'֟�L�s�>QΘ�z+54G���>�_�:�O��ª����G$��1��s�T!��0�0#A$�G_N5��&��T8����,��1�t��ž�O,�����(e���6팀��i�s���5���c�����e;k/�=����
���ЛE���B�Sy�D�q��X>��G�:n~�|�9� v��`'Pq�������iüd?